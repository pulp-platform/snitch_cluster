// Copyright 2020 ETH Zurich
    // SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
    //
    // Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
    // Florian Zaruba <zarubaf@iis.ee.ethz.ch>
    // Stefan Mach <smach@iis.ee.ethz.ch>
    // Thomas Benz <tbenz@iis.ee.ethz.ch>
    // Paul Scheffler <paulsc@iis.ee.ethz.ch>
    // Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
    //
    // AUTOMATICALLY GENERATED by gen_bootrom_param.py; edit the script instead.

    module bootrom #(
        parameter int unsigned AddrWidth = 32,
        parameter int unsigned DataWidth = 32,
        parameter int unsigned BootromSize = 65536
    )(
        input  logic                 clk_i,
        input  logic                 rst_ni,
        input  logic [AddrWidth-1:0] addr_i,
        output logic [DataWidth-1:0] data_o
    );
        logic [BootromSize-1:0][7:0] rom = '{
            {8'h00}, /* 0xffff */
            {8'h00}, /* 0xfffe */
            {8'h00}, /* 0xfffd */
            {8'h00}, /* 0xfffc */
            {8'h00}, /* 0xfffb */
            {8'h00}, /* 0xfffa */
            {8'h00}, /* 0xfff9 */
            {8'h00}, /* 0xfff8 */
            {8'h00}, /* 0xfff7 */
            {8'h00}, /* 0xfff6 */
            {8'h00}, /* 0xfff5 */
            {8'h00}, /* 0xfff4 */
            {8'h00}, /* 0xfff3 */
            {8'h00}, /* 0xfff2 */
            {8'h00}, /* 0xfff1 */
            {8'h00}, /* 0xfff0 */
            {8'h00}, /* 0xffef */
            {8'h00}, /* 0xffee */
            {8'h00}, /* 0xffed */
            {8'h00}, /* 0xffec */
            {8'h00}, /* 0xffeb */
            {8'h00}, /* 0xffea */
            {8'h00}, /* 0xffe9 */
            {8'h00}, /* 0xffe8 */
            {8'h00}, /* 0xffe7 */
            {8'h00}, /* 0xffe6 */
            {8'h00}, /* 0xffe5 */
            {8'h00}, /* 0xffe4 */
            {8'h00}, /* 0xffe3 */
            {8'h00}, /* 0xffe2 */
            {8'h00}, /* 0xffe1 */
            {8'h00}, /* 0xffe0 */
            {8'h00}, /* 0xffdf */
            {8'h00}, /* 0xffde */
            {8'h00}, /* 0xffdd */
            {8'h00}, /* 0xffdc */
            {8'h00}, /* 0xffdb */
            {8'h00}, /* 0xffda */
            {8'h00}, /* 0xffd9 */
            {8'h00}, /* 0xffd8 */
            {8'h00}, /* 0xffd7 */
            {8'h00}, /* 0xffd6 */
            {8'h00}, /* 0xffd5 */
            {8'h00}, /* 0xffd4 */
            {8'h00}, /* 0xffd3 */
            {8'h00}, /* 0xffd2 */
            {8'h00}, /* 0xffd1 */
            {8'h00}, /* 0xffd0 */
            {8'h00}, /* 0xffcf */
            {8'h00}, /* 0xffce */
            {8'h00}, /* 0xffcd */
            {8'h00}, /* 0xffcc */
            {8'h00}, /* 0xffcb */
            {8'h00}, /* 0xffca */
            {8'h00}, /* 0xffc9 */
            {8'h00}, /* 0xffc8 */
            {8'h00}, /* 0xffc7 */
            {8'h00}, /* 0xffc6 */
            {8'h00}, /* 0xffc5 */
            {8'h00}, /* 0xffc4 */
            {8'h00}, /* 0xffc3 */
            {8'h00}, /* 0xffc2 */
            {8'h00}, /* 0xffc1 */
            {8'h00}, /* 0xffc0 */
            {8'h00}, /* 0xffbf */
            {8'h00}, /* 0xffbe */
            {8'h00}, /* 0xffbd */
            {8'h00}, /* 0xffbc */
            {8'h00}, /* 0xffbb */
            {8'h00}, /* 0xffba */
            {8'h00}, /* 0xffb9 */
            {8'h00}, /* 0xffb8 */
            {8'h00}, /* 0xffb7 */
            {8'h00}, /* 0xffb6 */
            {8'h00}, /* 0xffb5 */
            {8'h00}, /* 0xffb4 */
            {8'h00}, /* 0xffb3 */
            {8'h00}, /* 0xffb2 */
            {8'h00}, /* 0xffb1 */
            {8'h00}, /* 0xffb0 */
            {8'h00}, /* 0xffaf */
            {8'h00}, /* 0xffae */
            {8'h00}, /* 0xffad */
            {8'h00}, /* 0xffac */
            {8'h00}, /* 0xffab */
            {8'h00}, /* 0xffaa */
            {8'h00}, /* 0xffa9 */
            {8'h00}, /* 0xffa8 */
            {8'h00}, /* 0xffa7 */
            {8'h00}, /* 0xffa6 */
            {8'h00}, /* 0xffa5 */
            {8'h00}, /* 0xffa4 */
            {8'h00}, /* 0xffa3 */
            {8'h00}, /* 0xffa2 */
            {8'h00}, /* 0xffa1 */
            {8'h00}, /* 0xffa0 */
            {8'h00}, /* 0xff9f */
            {8'h00}, /* 0xff9e */
            {8'h00}, /* 0xff9d */
            {8'h00}, /* 0xff9c */
            {8'h00}, /* 0xff9b */
            {8'h00}, /* 0xff9a */
            {8'h00}, /* 0xff99 */
            {8'h00}, /* 0xff98 */
            {8'h00}, /* 0xff97 */
            {8'h00}, /* 0xff96 */
            {8'h00}, /* 0xff95 */
            {8'h00}, /* 0xff94 */
            {8'h00}, /* 0xff93 */
            {8'h00}, /* 0xff92 */
            {8'h00}, /* 0xff91 */
            {8'h00}, /* 0xff90 */
            {8'h00}, /* 0xff8f */
            {8'h00}, /* 0xff8e */
            {8'h00}, /* 0xff8d */
            {8'h00}, /* 0xff8c */
            {8'h00}, /* 0xff8b */
            {8'h00}, /* 0xff8a */
            {8'h00}, /* 0xff89 */
            {8'h00}, /* 0xff88 */
            {8'h00}, /* 0xff87 */
            {8'h00}, /* 0xff86 */
            {8'h00}, /* 0xff85 */
            {8'h00}, /* 0xff84 */
            {8'h00}, /* 0xff83 */
            {8'h00}, /* 0xff82 */
            {8'h00}, /* 0xff81 */
            {8'h00}, /* 0xff80 */
            {8'h00}, /* 0xff7f */
            {8'h00}, /* 0xff7e */
            {8'h00}, /* 0xff7d */
            {8'h00}, /* 0xff7c */
            {8'h00}, /* 0xff7b */
            {8'h00}, /* 0xff7a */
            {8'h00}, /* 0xff79 */
            {8'h00}, /* 0xff78 */
            {8'h00}, /* 0xff77 */
            {8'h00}, /* 0xff76 */
            {8'h00}, /* 0xff75 */
            {8'h00}, /* 0xff74 */
            {8'h00}, /* 0xff73 */
            {8'h00}, /* 0xff72 */
            {8'h00}, /* 0xff71 */
            {8'h00}, /* 0xff70 */
            {8'h00}, /* 0xff6f */
            {8'h00}, /* 0xff6e */
            {8'h00}, /* 0xff6d */
            {8'h00}, /* 0xff6c */
            {8'h00}, /* 0xff6b */
            {8'h00}, /* 0xff6a */
            {8'h00}, /* 0xff69 */
            {8'h00}, /* 0xff68 */
            {8'h00}, /* 0xff67 */
            {8'h00}, /* 0xff66 */
            {8'h00}, /* 0xff65 */
            {8'h00}, /* 0xff64 */
            {8'h00}, /* 0xff63 */
            {8'h00}, /* 0xff62 */
            {8'h00}, /* 0xff61 */
            {8'h00}, /* 0xff60 */
            {8'h00}, /* 0xff5f */
            {8'h00}, /* 0xff5e */
            {8'h00}, /* 0xff5d */
            {8'h00}, /* 0xff5c */
            {8'h00}, /* 0xff5b */
            {8'h00}, /* 0xff5a */
            {8'h00}, /* 0xff59 */
            {8'h00}, /* 0xff58 */
            {8'h00}, /* 0xff57 */
            {8'h00}, /* 0xff56 */
            {8'h00}, /* 0xff55 */
            {8'h00}, /* 0xff54 */
            {8'h00}, /* 0xff53 */
            {8'h00}, /* 0xff52 */
            {8'h00}, /* 0xff51 */
            {8'h00}, /* 0xff50 */
            {8'h00}, /* 0xff4f */
            {8'h00}, /* 0xff4e */
            {8'h00}, /* 0xff4d */
            {8'h00}, /* 0xff4c */
            {8'h00}, /* 0xff4b */
            {8'h00}, /* 0xff4a */
            {8'h00}, /* 0xff49 */
            {8'h00}, /* 0xff48 */
            {8'h00}, /* 0xff47 */
            {8'h00}, /* 0xff46 */
            {8'h00}, /* 0xff45 */
            {8'h00}, /* 0xff44 */
            {8'h00}, /* 0xff43 */
            {8'h00}, /* 0xff42 */
            {8'h00}, /* 0xff41 */
            {8'h00}, /* 0xff40 */
            {8'h00}, /* 0xff3f */
            {8'h00}, /* 0xff3e */
            {8'h00}, /* 0xff3d */
            {8'h00}, /* 0xff3c */
            {8'h00}, /* 0xff3b */
            {8'h00}, /* 0xff3a */
            {8'h00}, /* 0xff39 */
            {8'h00}, /* 0xff38 */
            {8'h00}, /* 0xff37 */
            {8'h00}, /* 0xff36 */
            {8'h00}, /* 0xff35 */
            {8'h00}, /* 0xff34 */
            {8'h00}, /* 0xff33 */
            {8'h00}, /* 0xff32 */
            {8'h00}, /* 0xff31 */
            {8'h00}, /* 0xff30 */
            {8'h00}, /* 0xff2f */
            {8'h00}, /* 0xff2e */
            {8'h00}, /* 0xff2d */
            {8'h00}, /* 0xff2c */
            {8'h00}, /* 0xff2b */
            {8'h00}, /* 0xff2a */
            {8'h00}, /* 0xff29 */
            {8'h00}, /* 0xff28 */
            {8'h00}, /* 0xff27 */
            {8'h00}, /* 0xff26 */
            {8'h00}, /* 0xff25 */
            {8'h00}, /* 0xff24 */
            {8'h00}, /* 0xff23 */
            {8'h00}, /* 0xff22 */
            {8'h00}, /* 0xff21 */
            {8'h00}, /* 0xff20 */
            {8'h00}, /* 0xff1f */
            {8'h00}, /* 0xff1e */
            {8'h00}, /* 0xff1d */
            {8'h00}, /* 0xff1c */
            {8'h00}, /* 0xff1b */
            {8'h00}, /* 0xff1a */
            {8'h00}, /* 0xff19 */
            {8'h00}, /* 0xff18 */
            {8'h00}, /* 0xff17 */
            {8'h00}, /* 0xff16 */
            {8'h00}, /* 0xff15 */
            {8'h00}, /* 0xff14 */
            {8'h00}, /* 0xff13 */
            {8'h00}, /* 0xff12 */
            {8'h00}, /* 0xff11 */
            {8'h00}, /* 0xff10 */
            {8'h00}, /* 0xff0f */
            {8'h00}, /* 0xff0e */
            {8'h00}, /* 0xff0d */
            {8'h00}, /* 0xff0c */
            {8'h00}, /* 0xff0b */
            {8'h00}, /* 0xff0a */
            {8'h00}, /* 0xff09 */
            {8'h00}, /* 0xff08 */
            {8'h00}, /* 0xff07 */
            {8'h00}, /* 0xff06 */
            {8'h00}, /* 0xff05 */
            {8'h00}, /* 0xff04 */
            {8'h00}, /* 0xff03 */
            {8'h00}, /* 0xff02 */
            {8'h00}, /* 0xff01 */
            {8'h00}, /* 0xff00 */
            {8'h00}, /* 0xfeff */
            {8'h00}, /* 0xfefe */
            {8'h00}, /* 0xfefd */
            {8'h00}, /* 0xfefc */
            {8'h00}, /* 0xfefb */
            {8'h00}, /* 0xfefa */
            {8'h00}, /* 0xfef9 */
            {8'h00}, /* 0xfef8 */
            {8'h00}, /* 0xfef7 */
            {8'h00}, /* 0xfef6 */
            {8'h00}, /* 0xfef5 */
            {8'h00}, /* 0xfef4 */
            {8'h00}, /* 0xfef3 */
            {8'h00}, /* 0xfef2 */
            {8'h00}, /* 0xfef1 */
            {8'h00}, /* 0xfef0 */
            {8'h00}, /* 0xfeef */
            {8'h00}, /* 0xfeee */
            {8'h00}, /* 0xfeed */
            {8'h00}, /* 0xfeec */
            {8'h00}, /* 0xfeeb */
            {8'h00}, /* 0xfeea */
            {8'h00}, /* 0xfee9 */
            {8'h00}, /* 0xfee8 */
            {8'h00}, /* 0xfee7 */
            {8'h00}, /* 0xfee6 */
            {8'h00}, /* 0xfee5 */
            {8'h00}, /* 0xfee4 */
            {8'h00}, /* 0xfee3 */
            {8'h00}, /* 0xfee2 */
            {8'h00}, /* 0xfee1 */
            {8'h00}, /* 0xfee0 */
            {8'h00}, /* 0xfedf */
            {8'h00}, /* 0xfede */
            {8'h00}, /* 0xfedd */
            {8'h00}, /* 0xfedc */
            {8'h00}, /* 0xfedb */
            {8'h00}, /* 0xfeda */
            {8'h00}, /* 0xfed9 */
            {8'h00}, /* 0xfed8 */
            {8'h00}, /* 0xfed7 */
            {8'h00}, /* 0xfed6 */
            {8'h00}, /* 0xfed5 */
            {8'h00}, /* 0xfed4 */
            {8'h00}, /* 0xfed3 */
            {8'h00}, /* 0xfed2 */
            {8'h00}, /* 0xfed1 */
            {8'h00}, /* 0xfed0 */
            {8'h00}, /* 0xfecf */
            {8'h00}, /* 0xfece */
            {8'h00}, /* 0xfecd */
            {8'h00}, /* 0xfecc */
            {8'h00}, /* 0xfecb */
            {8'h00}, /* 0xfeca */
            {8'h00}, /* 0xfec9 */
            {8'h00}, /* 0xfec8 */
            {8'h00}, /* 0xfec7 */
            {8'h00}, /* 0xfec6 */
            {8'h00}, /* 0xfec5 */
            {8'h00}, /* 0xfec4 */
            {8'h00}, /* 0xfec3 */
            {8'h00}, /* 0xfec2 */
            {8'h00}, /* 0xfec1 */
            {8'h00}, /* 0xfec0 */
            {8'h00}, /* 0xfebf */
            {8'h00}, /* 0xfebe */
            {8'h00}, /* 0xfebd */
            {8'h00}, /* 0xfebc */
            {8'h00}, /* 0xfebb */
            {8'h00}, /* 0xfeba */
            {8'h00}, /* 0xfeb9 */
            {8'h00}, /* 0xfeb8 */
            {8'h00}, /* 0xfeb7 */
            {8'h00}, /* 0xfeb6 */
            {8'h00}, /* 0xfeb5 */
            {8'h00}, /* 0xfeb4 */
            {8'h00}, /* 0xfeb3 */
            {8'h00}, /* 0xfeb2 */
            {8'h00}, /* 0xfeb1 */
            {8'h00}, /* 0xfeb0 */
            {8'h00}, /* 0xfeaf */
            {8'h00}, /* 0xfeae */
            {8'h00}, /* 0xfead */
            {8'h00}, /* 0xfeac */
            {8'h00}, /* 0xfeab */
            {8'h00}, /* 0xfeaa */
            {8'h00}, /* 0xfea9 */
            {8'h00}, /* 0xfea8 */
            {8'h00}, /* 0xfea7 */
            {8'h00}, /* 0xfea6 */
            {8'h00}, /* 0xfea5 */
            {8'h00}, /* 0xfea4 */
            {8'h00}, /* 0xfea3 */
            {8'h00}, /* 0xfea2 */
            {8'h00}, /* 0xfea1 */
            {8'h00}, /* 0xfea0 */
            {8'h00}, /* 0xfe9f */
            {8'h00}, /* 0xfe9e */
            {8'h00}, /* 0xfe9d */
            {8'h00}, /* 0xfe9c */
            {8'h00}, /* 0xfe9b */
            {8'h00}, /* 0xfe9a */
            {8'h00}, /* 0xfe99 */
            {8'h00}, /* 0xfe98 */
            {8'h00}, /* 0xfe97 */
            {8'h00}, /* 0xfe96 */
            {8'h00}, /* 0xfe95 */
            {8'h00}, /* 0xfe94 */
            {8'h00}, /* 0xfe93 */
            {8'h00}, /* 0xfe92 */
            {8'h00}, /* 0xfe91 */
            {8'h00}, /* 0xfe90 */
            {8'h00}, /* 0xfe8f */
            {8'h00}, /* 0xfe8e */
            {8'h00}, /* 0xfe8d */
            {8'h00}, /* 0xfe8c */
            {8'h00}, /* 0xfe8b */
            {8'h00}, /* 0xfe8a */
            {8'h00}, /* 0xfe89 */
            {8'h00}, /* 0xfe88 */
            {8'h00}, /* 0xfe87 */
            {8'h00}, /* 0xfe86 */
            {8'h00}, /* 0xfe85 */
            {8'h00}, /* 0xfe84 */
            {8'h00}, /* 0xfe83 */
            {8'h00}, /* 0xfe82 */
            {8'h00}, /* 0xfe81 */
            {8'h00}, /* 0xfe80 */
            {8'h00}, /* 0xfe7f */
            {8'h00}, /* 0xfe7e */
            {8'h00}, /* 0xfe7d */
            {8'h00}, /* 0xfe7c */
            {8'h00}, /* 0xfe7b */
            {8'h00}, /* 0xfe7a */
            {8'h00}, /* 0xfe79 */
            {8'h00}, /* 0xfe78 */
            {8'h00}, /* 0xfe77 */
            {8'h00}, /* 0xfe76 */
            {8'h00}, /* 0xfe75 */
            {8'h00}, /* 0xfe74 */
            {8'h00}, /* 0xfe73 */
            {8'h00}, /* 0xfe72 */
            {8'h00}, /* 0xfe71 */
            {8'h00}, /* 0xfe70 */
            {8'h00}, /* 0xfe6f */
            {8'h00}, /* 0xfe6e */
            {8'h00}, /* 0xfe6d */
            {8'h00}, /* 0xfe6c */
            {8'h00}, /* 0xfe6b */
            {8'h00}, /* 0xfe6a */
            {8'h00}, /* 0xfe69 */
            {8'h00}, /* 0xfe68 */
            {8'h00}, /* 0xfe67 */
            {8'h00}, /* 0xfe66 */
            {8'h00}, /* 0xfe65 */
            {8'h00}, /* 0xfe64 */
            {8'h00}, /* 0xfe63 */
            {8'h00}, /* 0xfe62 */
            {8'h00}, /* 0xfe61 */
            {8'h00}, /* 0xfe60 */
            {8'h00}, /* 0xfe5f */
            {8'h00}, /* 0xfe5e */
            {8'h00}, /* 0xfe5d */
            {8'h00}, /* 0xfe5c */
            {8'h00}, /* 0xfe5b */
            {8'h00}, /* 0xfe5a */
            {8'h00}, /* 0xfe59 */
            {8'h00}, /* 0xfe58 */
            {8'h00}, /* 0xfe57 */
            {8'h00}, /* 0xfe56 */
            {8'h00}, /* 0xfe55 */
            {8'h00}, /* 0xfe54 */
            {8'h00}, /* 0xfe53 */
            {8'h00}, /* 0xfe52 */
            {8'h00}, /* 0xfe51 */
            {8'h00}, /* 0xfe50 */
            {8'h00}, /* 0xfe4f */
            {8'h00}, /* 0xfe4e */
            {8'h00}, /* 0xfe4d */
            {8'h00}, /* 0xfe4c */
            {8'h00}, /* 0xfe4b */
            {8'h00}, /* 0xfe4a */
            {8'h00}, /* 0xfe49 */
            {8'h00}, /* 0xfe48 */
            {8'h00}, /* 0xfe47 */
            {8'h00}, /* 0xfe46 */
            {8'h00}, /* 0xfe45 */
            {8'h00}, /* 0xfe44 */
            {8'h00}, /* 0xfe43 */
            {8'h00}, /* 0xfe42 */
            {8'h00}, /* 0xfe41 */
            {8'h00}, /* 0xfe40 */
            {8'h00}, /* 0xfe3f */
            {8'h00}, /* 0xfe3e */
            {8'h00}, /* 0xfe3d */
            {8'h00}, /* 0xfe3c */
            {8'h00}, /* 0xfe3b */
            {8'h00}, /* 0xfe3a */
            {8'h00}, /* 0xfe39 */
            {8'h00}, /* 0xfe38 */
            {8'h00}, /* 0xfe37 */
            {8'h00}, /* 0xfe36 */
            {8'h00}, /* 0xfe35 */
            {8'h00}, /* 0xfe34 */
            {8'h00}, /* 0xfe33 */
            {8'h00}, /* 0xfe32 */
            {8'h00}, /* 0xfe31 */
            {8'h00}, /* 0xfe30 */
            {8'h00}, /* 0xfe2f */
            {8'h00}, /* 0xfe2e */
            {8'h00}, /* 0xfe2d */
            {8'h00}, /* 0xfe2c */
            {8'h00}, /* 0xfe2b */
            {8'h00}, /* 0xfe2a */
            {8'h00}, /* 0xfe29 */
            {8'h00}, /* 0xfe28 */
            {8'h00}, /* 0xfe27 */
            {8'h00}, /* 0xfe26 */
            {8'h00}, /* 0xfe25 */
            {8'h00}, /* 0xfe24 */
            {8'h00}, /* 0xfe23 */
            {8'h00}, /* 0xfe22 */
            {8'h00}, /* 0xfe21 */
            {8'h00}, /* 0xfe20 */
            {8'h00}, /* 0xfe1f */
            {8'h00}, /* 0xfe1e */
            {8'h00}, /* 0xfe1d */
            {8'h00}, /* 0xfe1c */
            {8'h00}, /* 0xfe1b */
            {8'h00}, /* 0xfe1a */
            {8'h00}, /* 0xfe19 */
            {8'h00}, /* 0xfe18 */
            {8'h00}, /* 0xfe17 */
            {8'h00}, /* 0xfe16 */
            {8'h00}, /* 0xfe15 */
            {8'h00}, /* 0xfe14 */
            {8'h00}, /* 0xfe13 */
            {8'h00}, /* 0xfe12 */
            {8'h00}, /* 0xfe11 */
            {8'h00}, /* 0xfe10 */
            {8'h00}, /* 0xfe0f */
            {8'h00}, /* 0xfe0e */
            {8'h00}, /* 0xfe0d */
            {8'h00}, /* 0xfe0c */
            {8'h00}, /* 0xfe0b */
            {8'h00}, /* 0xfe0a */
            {8'h00}, /* 0xfe09 */
            {8'h00}, /* 0xfe08 */
            {8'h00}, /* 0xfe07 */
            {8'h00}, /* 0xfe06 */
            {8'h00}, /* 0xfe05 */
            {8'h00}, /* 0xfe04 */
            {8'h00}, /* 0xfe03 */
            {8'h00}, /* 0xfe02 */
            {8'h00}, /* 0xfe01 */
            {8'h00}, /* 0xfe00 */
            {8'h00}, /* 0xfdff */
            {8'h00}, /* 0xfdfe */
            {8'h00}, /* 0xfdfd */
            {8'h00}, /* 0xfdfc */
            {8'h00}, /* 0xfdfb */
            {8'h00}, /* 0xfdfa */
            {8'h00}, /* 0xfdf9 */
            {8'h00}, /* 0xfdf8 */
            {8'h00}, /* 0xfdf7 */
            {8'h00}, /* 0xfdf6 */
            {8'h00}, /* 0xfdf5 */
            {8'h00}, /* 0xfdf4 */
            {8'h00}, /* 0xfdf3 */
            {8'h00}, /* 0xfdf2 */
            {8'h00}, /* 0xfdf1 */
            {8'h00}, /* 0xfdf0 */
            {8'h00}, /* 0xfdef */
            {8'h00}, /* 0xfdee */
            {8'h00}, /* 0xfded */
            {8'h00}, /* 0xfdec */
            {8'h00}, /* 0xfdeb */
            {8'h00}, /* 0xfdea */
            {8'h00}, /* 0xfde9 */
            {8'h00}, /* 0xfde8 */
            {8'h00}, /* 0xfde7 */
            {8'h00}, /* 0xfde6 */
            {8'h00}, /* 0xfde5 */
            {8'h00}, /* 0xfde4 */
            {8'h00}, /* 0xfde3 */
            {8'h00}, /* 0xfde2 */
            {8'h00}, /* 0xfde1 */
            {8'h00}, /* 0xfde0 */
            {8'h00}, /* 0xfddf */
            {8'h00}, /* 0xfdde */
            {8'h00}, /* 0xfddd */
            {8'h00}, /* 0xfddc */
            {8'h00}, /* 0xfddb */
            {8'h00}, /* 0xfdda */
            {8'h00}, /* 0xfdd9 */
            {8'h00}, /* 0xfdd8 */
            {8'h00}, /* 0xfdd7 */
            {8'h00}, /* 0xfdd6 */
            {8'h00}, /* 0xfdd5 */
            {8'h00}, /* 0xfdd4 */
            {8'h00}, /* 0xfdd3 */
            {8'h00}, /* 0xfdd2 */
            {8'h00}, /* 0xfdd1 */
            {8'h00}, /* 0xfdd0 */
            {8'h00}, /* 0xfdcf */
            {8'h00}, /* 0xfdce */
            {8'h00}, /* 0xfdcd */
            {8'h00}, /* 0xfdcc */
            {8'h00}, /* 0xfdcb */
            {8'h00}, /* 0xfdca */
            {8'h00}, /* 0xfdc9 */
            {8'h00}, /* 0xfdc8 */
            {8'h00}, /* 0xfdc7 */
            {8'h00}, /* 0xfdc6 */
            {8'h00}, /* 0xfdc5 */
            {8'h00}, /* 0xfdc4 */
            {8'h00}, /* 0xfdc3 */
            {8'h00}, /* 0xfdc2 */
            {8'h00}, /* 0xfdc1 */
            {8'h00}, /* 0xfdc0 */
            {8'h00}, /* 0xfdbf */
            {8'h00}, /* 0xfdbe */
            {8'h00}, /* 0xfdbd */
            {8'h00}, /* 0xfdbc */
            {8'h00}, /* 0xfdbb */
            {8'h00}, /* 0xfdba */
            {8'h00}, /* 0xfdb9 */
            {8'h00}, /* 0xfdb8 */
            {8'h00}, /* 0xfdb7 */
            {8'h00}, /* 0xfdb6 */
            {8'h00}, /* 0xfdb5 */
            {8'h00}, /* 0xfdb4 */
            {8'h00}, /* 0xfdb3 */
            {8'h00}, /* 0xfdb2 */
            {8'h00}, /* 0xfdb1 */
            {8'h00}, /* 0xfdb0 */
            {8'h00}, /* 0xfdaf */
            {8'h00}, /* 0xfdae */
            {8'h00}, /* 0xfdad */
            {8'h00}, /* 0xfdac */
            {8'h00}, /* 0xfdab */
            {8'h00}, /* 0xfdaa */
            {8'h00}, /* 0xfda9 */
            {8'h00}, /* 0xfda8 */
            {8'h00}, /* 0xfda7 */
            {8'h00}, /* 0xfda6 */
            {8'h00}, /* 0xfda5 */
            {8'h00}, /* 0xfda4 */
            {8'h00}, /* 0xfda3 */
            {8'h00}, /* 0xfda2 */
            {8'h00}, /* 0xfda1 */
            {8'h00}, /* 0xfda0 */
            {8'h00}, /* 0xfd9f */
            {8'h00}, /* 0xfd9e */
            {8'h00}, /* 0xfd9d */
            {8'h00}, /* 0xfd9c */
            {8'h00}, /* 0xfd9b */
            {8'h00}, /* 0xfd9a */
            {8'h00}, /* 0xfd99 */
            {8'h00}, /* 0xfd98 */
            {8'h00}, /* 0xfd97 */
            {8'h00}, /* 0xfd96 */
            {8'h00}, /* 0xfd95 */
            {8'h00}, /* 0xfd94 */
            {8'h00}, /* 0xfd93 */
            {8'h00}, /* 0xfd92 */
            {8'h00}, /* 0xfd91 */
            {8'h00}, /* 0xfd90 */
            {8'h00}, /* 0xfd8f */
            {8'h00}, /* 0xfd8e */
            {8'h00}, /* 0xfd8d */
            {8'h00}, /* 0xfd8c */
            {8'h00}, /* 0xfd8b */
            {8'h00}, /* 0xfd8a */
            {8'h00}, /* 0xfd89 */
            {8'h00}, /* 0xfd88 */
            {8'h00}, /* 0xfd87 */
            {8'h00}, /* 0xfd86 */
            {8'h00}, /* 0xfd85 */
            {8'h00}, /* 0xfd84 */
            {8'h00}, /* 0xfd83 */
            {8'h00}, /* 0xfd82 */
            {8'h00}, /* 0xfd81 */
            {8'h00}, /* 0xfd80 */
            {8'h00}, /* 0xfd7f */
            {8'h00}, /* 0xfd7e */
            {8'h00}, /* 0xfd7d */
            {8'h00}, /* 0xfd7c */
            {8'h00}, /* 0xfd7b */
            {8'h00}, /* 0xfd7a */
            {8'h00}, /* 0xfd79 */
            {8'h00}, /* 0xfd78 */
            {8'h00}, /* 0xfd77 */
            {8'h00}, /* 0xfd76 */
            {8'h00}, /* 0xfd75 */
            {8'h00}, /* 0xfd74 */
            {8'h00}, /* 0xfd73 */
            {8'h00}, /* 0xfd72 */
            {8'h00}, /* 0xfd71 */
            {8'h00}, /* 0xfd70 */
            {8'h00}, /* 0xfd6f */
            {8'h00}, /* 0xfd6e */
            {8'h00}, /* 0xfd6d */
            {8'h00}, /* 0xfd6c */
            {8'h00}, /* 0xfd6b */
            {8'h00}, /* 0xfd6a */
            {8'h00}, /* 0xfd69 */
            {8'h00}, /* 0xfd68 */
            {8'h00}, /* 0xfd67 */
            {8'h00}, /* 0xfd66 */
            {8'h00}, /* 0xfd65 */
            {8'h00}, /* 0xfd64 */
            {8'h00}, /* 0xfd63 */
            {8'h00}, /* 0xfd62 */
            {8'h00}, /* 0xfd61 */
            {8'h00}, /* 0xfd60 */
            {8'h00}, /* 0xfd5f */
            {8'h00}, /* 0xfd5e */
            {8'h00}, /* 0xfd5d */
            {8'h00}, /* 0xfd5c */
            {8'h00}, /* 0xfd5b */
            {8'h00}, /* 0xfd5a */
            {8'h00}, /* 0xfd59 */
            {8'h00}, /* 0xfd58 */
            {8'h00}, /* 0xfd57 */
            {8'h00}, /* 0xfd56 */
            {8'h00}, /* 0xfd55 */
            {8'h00}, /* 0xfd54 */
            {8'h00}, /* 0xfd53 */
            {8'h00}, /* 0xfd52 */
            {8'h00}, /* 0xfd51 */
            {8'h00}, /* 0xfd50 */
            {8'h00}, /* 0xfd4f */
            {8'h00}, /* 0xfd4e */
            {8'h00}, /* 0xfd4d */
            {8'h00}, /* 0xfd4c */
            {8'h00}, /* 0xfd4b */
            {8'h00}, /* 0xfd4a */
            {8'h00}, /* 0xfd49 */
            {8'h00}, /* 0xfd48 */
            {8'h00}, /* 0xfd47 */
            {8'h00}, /* 0xfd46 */
            {8'h00}, /* 0xfd45 */
            {8'h00}, /* 0xfd44 */
            {8'h00}, /* 0xfd43 */
            {8'h00}, /* 0xfd42 */
            {8'h00}, /* 0xfd41 */
            {8'h00}, /* 0xfd40 */
            {8'h00}, /* 0xfd3f */
            {8'h00}, /* 0xfd3e */
            {8'h00}, /* 0xfd3d */
            {8'h00}, /* 0xfd3c */
            {8'h00}, /* 0xfd3b */
            {8'h00}, /* 0xfd3a */
            {8'h00}, /* 0xfd39 */
            {8'h00}, /* 0xfd38 */
            {8'h00}, /* 0xfd37 */
            {8'h00}, /* 0xfd36 */
            {8'h00}, /* 0xfd35 */
            {8'h00}, /* 0xfd34 */
            {8'h00}, /* 0xfd33 */
            {8'h00}, /* 0xfd32 */
            {8'h00}, /* 0xfd31 */
            {8'h00}, /* 0xfd30 */
            {8'h00}, /* 0xfd2f */
            {8'h00}, /* 0xfd2e */
            {8'h00}, /* 0xfd2d */
            {8'h00}, /* 0xfd2c */
            {8'h00}, /* 0xfd2b */
            {8'h00}, /* 0xfd2a */
            {8'h00}, /* 0xfd29 */
            {8'h00}, /* 0xfd28 */
            {8'h00}, /* 0xfd27 */
            {8'h00}, /* 0xfd26 */
            {8'h00}, /* 0xfd25 */
            {8'h00}, /* 0xfd24 */
            {8'h00}, /* 0xfd23 */
            {8'h00}, /* 0xfd22 */
            {8'h00}, /* 0xfd21 */
            {8'h00}, /* 0xfd20 */
            {8'h00}, /* 0xfd1f */
            {8'h00}, /* 0xfd1e */
            {8'h00}, /* 0xfd1d */
            {8'h00}, /* 0xfd1c */
            {8'h00}, /* 0xfd1b */
            {8'h00}, /* 0xfd1a */
            {8'h00}, /* 0xfd19 */
            {8'h00}, /* 0xfd18 */
            {8'h00}, /* 0xfd17 */
            {8'h00}, /* 0xfd16 */
            {8'h00}, /* 0xfd15 */
            {8'h00}, /* 0xfd14 */
            {8'h00}, /* 0xfd13 */
            {8'h00}, /* 0xfd12 */
            {8'h00}, /* 0xfd11 */
            {8'h00}, /* 0xfd10 */
            {8'h00}, /* 0xfd0f */
            {8'h00}, /* 0xfd0e */
            {8'h00}, /* 0xfd0d */
            {8'h00}, /* 0xfd0c */
            {8'h00}, /* 0xfd0b */
            {8'h00}, /* 0xfd0a */
            {8'h00}, /* 0xfd09 */
            {8'h00}, /* 0xfd08 */
            {8'h00}, /* 0xfd07 */
            {8'h00}, /* 0xfd06 */
            {8'h00}, /* 0xfd05 */
            {8'h00}, /* 0xfd04 */
            {8'h00}, /* 0xfd03 */
            {8'h00}, /* 0xfd02 */
            {8'h00}, /* 0xfd01 */
            {8'h00}, /* 0xfd00 */
            {8'h00}, /* 0xfcff */
            {8'h00}, /* 0xfcfe */
            {8'h00}, /* 0xfcfd */
            {8'h00}, /* 0xfcfc */
            {8'h00}, /* 0xfcfb */
            {8'h00}, /* 0xfcfa */
            {8'h00}, /* 0xfcf9 */
            {8'h00}, /* 0xfcf8 */
            {8'h00}, /* 0xfcf7 */
            {8'h00}, /* 0xfcf6 */
            {8'h00}, /* 0xfcf5 */
            {8'h00}, /* 0xfcf4 */
            {8'h00}, /* 0xfcf3 */
            {8'h00}, /* 0xfcf2 */
            {8'h00}, /* 0xfcf1 */
            {8'h00}, /* 0xfcf0 */
            {8'h00}, /* 0xfcef */
            {8'h00}, /* 0xfcee */
            {8'h00}, /* 0xfced */
            {8'h00}, /* 0xfcec */
            {8'h00}, /* 0xfceb */
            {8'h00}, /* 0xfcea */
            {8'h00}, /* 0xfce9 */
            {8'h00}, /* 0xfce8 */
            {8'h00}, /* 0xfce7 */
            {8'h00}, /* 0xfce6 */
            {8'h00}, /* 0xfce5 */
            {8'h00}, /* 0xfce4 */
            {8'h00}, /* 0xfce3 */
            {8'h00}, /* 0xfce2 */
            {8'h00}, /* 0xfce1 */
            {8'h00}, /* 0xfce0 */
            {8'h00}, /* 0xfcdf */
            {8'h00}, /* 0xfcde */
            {8'h00}, /* 0xfcdd */
            {8'h00}, /* 0xfcdc */
            {8'h00}, /* 0xfcdb */
            {8'h00}, /* 0xfcda */
            {8'h00}, /* 0xfcd9 */
            {8'h00}, /* 0xfcd8 */
            {8'h00}, /* 0xfcd7 */
            {8'h00}, /* 0xfcd6 */
            {8'h00}, /* 0xfcd5 */
            {8'h00}, /* 0xfcd4 */
            {8'h00}, /* 0xfcd3 */
            {8'h00}, /* 0xfcd2 */
            {8'h00}, /* 0xfcd1 */
            {8'h00}, /* 0xfcd0 */
            {8'h00}, /* 0xfccf */
            {8'h00}, /* 0xfcce */
            {8'h00}, /* 0xfccd */
            {8'h00}, /* 0xfccc */
            {8'h00}, /* 0xfccb */
            {8'h00}, /* 0xfcca */
            {8'h00}, /* 0xfcc9 */
            {8'h00}, /* 0xfcc8 */
            {8'h00}, /* 0xfcc7 */
            {8'h00}, /* 0xfcc6 */
            {8'h00}, /* 0xfcc5 */
            {8'h00}, /* 0xfcc4 */
            {8'h00}, /* 0xfcc3 */
            {8'h00}, /* 0xfcc2 */
            {8'h00}, /* 0xfcc1 */
            {8'h00}, /* 0xfcc0 */
            {8'h00}, /* 0xfcbf */
            {8'h00}, /* 0xfcbe */
            {8'h00}, /* 0xfcbd */
            {8'h00}, /* 0xfcbc */
            {8'h00}, /* 0xfcbb */
            {8'h00}, /* 0xfcba */
            {8'h00}, /* 0xfcb9 */
            {8'h00}, /* 0xfcb8 */
            {8'h00}, /* 0xfcb7 */
            {8'h00}, /* 0xfcb6 */
            {8'h00}, /* 0xfcb5 */
            {8'h00}, /* 0xfcb4 */
            {8'h00}, /* 0xfcb3 */
            {8'h00}, /* 0xfcb2 */
            {8'h00}, /* 0xfcb1 */
            {8'h00}, /* 0xfcb0 */
            {8'h00}, /* 0xfcaf */
            {8'h00}, /* 0xfcae */
            {8'h00}, /* 0xfcad */
            {8'h00}, /* 0xfcac */
            {8'h00}, /* 0xfcab */
            {8'h00}, /* 0xfcaa */
            {8'h00}, /* 0xfca9 */
            {8'h00}, /* 0xfca8 */
            {8'h00}, /* 0xfca7 */
            {8'h00}, /* 0xfca6 */
            {8'h00}, /* 0xfca5 */
            {8'h00}, /* 0xfca4 */
            {8'h00}, /* 0xfca3 */
            {8'h00}, /* 0xfca2 */
            {8'h00}, /* 0xfca1 */
            {8'h00}, /* 0xfca0 */
            {8'h00}, /* 0xfc9f */
            {8'h00}, /* 0xfc9e */
            {8'h00}, /* 0xfc9d */
            {8'h00}, /* 0xfc9c */
            {8'h00}, /* 0xfc9b */
            {8'h00}, /* 0xfc9a */
            {8'h00}, /* 0xfc99 */
            {8'h00}, /* 0xfc98 */
            {8'h00}, /* 0xfc97 */
            {8'h00}, /* 0xfc96 */
            {8'h00}, /* 0xfc95 */
            {8'h00}, /* 0xfc94 */
            {8'h00}, /* 0xfc93 */
            {8'h00}, /* 0xfc92 */
            {8'h00}, /* 0xfc91 */
            {8'h00}, /* 0xfc90 */
            {8'h00}, /* 0xfc8f */
            {8'h00}, /* 0xfc8e */
            {8'h00}, /* 0xfc8d */
            {8'h00}, /* 0xfc8c */
            {8'h00}, /* 0xfc8b */
            {8'h00}, /* 0xfc8a */
            {8'h00}, /* 0xfc89 */
            {8'h00}, /* 0xfc88 */
            {8'h00}, /* 0xfc87 */
            {8'h00}, /* 0xfc86 */
            {8'h00}, /* 0xfc85 */
            {8'h00}, /* 0xfc84 */
            {8'h00}, /* 0xfc83 */
            {8'h00}, /* 0xfc82 */
            {8'h00}, /* 0xfc81 */
            {8'h00}, /* 0xfc80 */
            {8'h00}, /* 0xfc7f */
            {8'h00}, /* 0xfc7e */
            {8'h00}, /* 0xfc7d */
            {8'h00}, /* 0xfc7c */
            {8'h00}, /* 0xfc7b */
            {8'h00}, /* 0xfc7a */
            {8'h00}, /* 0xfc79 */
            {8'h00}, /* 0xfc78 */
            {8'h00}, /* 0xfc77 */
            {8'h00}, /* 0xfc76 */
            {8'h00}, /* 0xfc75 */
            {8'h00}, /* 0xfc74 */
            {8'h00}, /* 0xfc73 */
            {8'h00}, /* 0xfc72 */
            {8'h00}, /* 0xfc71 */
            {8'h00}, /* 0xfc70 */
            {8'h00}, /* 0xfc6f */
            {8'h00}, /* 0xfc6e */
            {8'h00}, /* 0xfc6d */
            {8'h00}, /* 0xfc6c */
            {8'h00}, /* 0xfc6b */
            {8'h00}, /* 0xfc6a */
            {8'h00}, /* 0xfc69 */
            {8'h00}, /* 0xfc68 */
            {8'h00}, /* 0xfc67 */
            {8'h00}, /* 0xfc66 */
            {8'h00}, /* 0xfc65 */
            {8'h00}, /* 0xfc64 */
            {8'h00}, /* 0xfc63 */
            {8'h00}, /* 0xfc62 */
            {8'h00}, /* 0xfc61 */
            {8'h00}, /* 0xfc60 */
            {8'h00}, /* 0xfc5f */
            {8'h00}, /* 0xfc5e */
            {8'h00}, /* 0xfc5d */
            {8'h00}, /* 0xfc5c */
            {8'h00}, /* 0xfc5b */
            {8'h00}, /* 0xfc5a */
            {8'h00}, /* 0xfc59 */
            {8'h00}, /* 0xfc58 */
            {8'h00}, /* 0xfc57 */
            {8'h00}, /* 0xfc56 */
            {8'h00}, /* 0xfc55 */
            {8'h00}, /* 0xfc54 */
            {8'h00}, /* 0xfc53 */
            {8'h00}, /* 0xfc52 */
            {8'h00}, /* 0xfc51 */
            {8'h00}, /* 0xfc50 */
            {8'h00}, /* 0xfc4f */
            {8'h00}, /* 0xfc4e */
            {8'h00}, /* 0xfc4d */
            {8'h00}, /* 0xfc4c */
            {8'h00}, /* 0xfc4b */
            {8'h00}, /* 0xfc4a */
            {8'h00}, /* 0xfc49 */
            {8'h00}, /* 0xfc48 */
            {8'h00}, /* 0xfc47 */
            {8'h00}, /* 0xfc46 */
            {8'h00}, /* 0xfc45 */
            {8'h00}, /* 0xfc44 */
            {8'h00}, /* 0xfc43 */
            {8'h00}, /* 0xfc42 */
            {8'h00}, /* 0xfc41 */
            {8'h00}, /* 0xfc40 */
            {8'h00}, /* 0xfc3f */
            {8'h00}, /* 0xfc3e */
            {8'h00}, /* 0xfc3d */
            {8'h00}, /* 0xfc3c */
            {8'h00}, /* 0xfc3b */
            {8'h00}, /* 0xfc3a */
            {8'h00}, /* 0xfc39 */
            {8'h00}, /* 0xfc38 */
            {8'h00}, /* 0xfc37 */
            {8'h00}, /* 0xfc36 */
            {8'h00}, /* 0xfc35 */
            {8'h00}, /* 0xfc34 */
            {8'h00}, /* 0xfc33 */
            {8'h00}, /* 0xfc32 */
            {8'h00}, /* 0xfc31 */
            {8'h00}, /* 0xfc30 */
            {8'h00}, /* 0xfc2f */
            {8'h00}, /* 0xfc2e */
            {8'h00}, /* 0xfc2d */
            {8'h00}, /* 0xfc2c */
            {8'h00}, /* 0xfc2b */
            {8'h00}, /* 0xfc2a */
            {8'h00}, /* 0xfc29 */
            {8'h00}, /* 0xfc28 */
            {8'h00}, /* 0xfc27 */
            {8'h00}, /* 0xfc26 */
            {8'h00}, /* 0xfc25 */
            {8'h00}, /* 0xfc24 */
            {8'h00}, /* 0xfc23 */
            {8'h00}, /* 0xfc22 */
            {8'h00}, /* 0xfc21 */
            {8'h00}, /* 0xfc20 */
            {8'h00}, /* 0xfc1f */
            {8'h00}, /* 0xfc1e */
            {8'h00}, /* 0xfc1d */
            {8'h00}, /* 0xfc1c */
            {8'h00}, /* 0xfc1b */
            {8'h00}, /* 0xfc1a */
            {8'h00}, /* 0xfc19 */
            {8'h00}, /* 0xfc18 */
            {8'h00}, /* 0xfc17 */
            {8'h00}, /* 0xfc16 */
            {8'h00}, /* 0xfc15 */
            {8'h00}, /* 0xfc14 */
            {8'h00}, /* 0xfc13 */
            {8'h00}, /* 0xfc12 */
            {8'h00}, /* 0xfc11 */
            {8'h00}, /* 0xfc10 */
            {8'h00}, /* 0xfc0f */
            {8'h00}, /* 0xfc0e */
            {8'h00}, /* 0xfc0d */
            {8'h00}, /* 0xfc0c */
            {8'h00}, /* 0xfc0b */
            {8'h00}, /* 0xfc0a */
            {8'h00}, /* 0xfc09 */
            {8'h00}, /* 0xfc08 */
            {8'h00}, /* 0xfc07 */
            {8'h00}, /* 0xfc06 */
            {8'h00}, /* 0xfc05 */
            {8'h00}, /* 0xfc04 */
            {8'h00}, /* 0xfc03 */
            {8'h00}, /* 0xfc02 */
            {8'h00}, /* 0xfc01 */
            {8'h00}, /* 0xfc00 */
            {8'h00}, /* 0xfbff */
            {8'h00}, /* 0xfbfe */
            {8'h00}, /* 0xfbfd */
            {8'h00}, /* 0xfbfc */
            {8'h00}, /* 0xfbfb */
            {8'h00}, /* 0xfbfa */
            {8'h00}, /* 0xfbf9 */
            {8'h00}, /* 0xfbf8 */
            {8'h00}, /* 0xfbf7 */
            {8'h00}, /* 0xfbf6 */
            {8'h00}, /* 0xfbf5 */
            {8'h00}, /* 0xfbf4 */
            {8'h00}, /* 0xfbf3 */
            {8'h00}, /* 0xfbf2 */
            {8'h00}, /* 0xfbf1 */
            {8'h00}, /* 0xfbf0 */
            {8'h00}, /* 0xfbef */
            {8'h00}, /* 0xfbee */
            {8'h00}, /* 0xfbed */
            {8'h00}, /* 0xfbec */
            {8'h00}, /* 0xfbeb */
            {8'h00}, /* 0xfbea */
            {8'h00}, /* 0xfbe9 */
            {8'h00}, /* 0xfbe8 */
            {8'h00}, /* 0xfbe7 */
            {8'h00}, /* 0xfbe6 */
            {8'h00}, /* 0xfbe5 */
            {8'h00}, /* 0xfbe4 */
            {8'h00}, /* 0xfbe3 */
            {8'h00}, /* 0xfbe2 */
            {8'h00}, /* 0xfbe1 */
            {8'h00}, /* 0xfbe0 */
            {8'h00}, /* 0xfbdf */
            {8'h00}, /* 0xfbde */
            {8'h00}, /* 0xfbdd */
            {8'h00}, /* 0xfbdc */
            {8'h00}, /* 0xfbdb */
            {8'h00}, /* 0xfbda */
            {8'h00}, /* 0xfbd9 */
            {8'h00}, /* 0xfbd8 */
            {8'h00}, /* 0xfbd7 */
            {8'h00}, /* 0xfbd6 */
            {8'h00}, /* 0xfbd5 */
            {8'h00}, /* 0xfbd4 */
            {8'h00}, /* 0xfbd3 */
            {8'h00}, /* 0xfbd2 */
            {8'h00}, /* 0xfbd1 */
            {8'h00}, /* 0xfbd0 */
            {8'h00}, /* 0xfbcf */
            {8'h00}, /* 0xfbce */
            {8'h00}, /* 0xfbcd */
            {8'h00}, /* 0xfbcc */
            {8'h00}, /* 0xfbcb */
            {8'h00}, /* 0xfbca */
            {8'h00}, /* 0xfbc9 */
            {8'h00}, /* 0xfbc8 */
            {8'h00}, /* 0xfbc7 */
            {8'h00}, /* 0xfbc6 */
            {8'h00}, /* 0xfbc5 */
            {8'h00}, /* 0xfbc4 */
            {8'h00}, /* 0xfbc3 */
            {8'h00}, /* 0xfbc2 */
            {8'h00}, /* 0xfbc1 */
            {8'h00}, /* 0xfbc0 */
            {8'h00}, /* 0xfbbf */
            {8'h00}, /* 0xfbbe */
            {8'h00}, /* 0xfbbd */
            {8'h00}, /* 0xfbbc */
            {8'h00}, /* 0xfbbb */
            {8'h00}, /* 0xfbba */
            {8'h00}, /* 0xfbb9 */
            {8'h00}, /* 0xfbb8 */
            {8'h00}, /* 0xfbb7 */
            {8'h00}, /* 0xfbb6 */
            {8'h00}, /* 0xfbb5 */
            {8'h00}, /* 0xfbb4 */
            {8'h00}, /* 0xfbb3 */
            {8'h00}, /* 0xfbb2 */
            {8'h00}, /* 0xfbb1 */
            {8'h00}, /* 0xfbb0 */
            {8'h00}, /* 0xfbaf */
            {8'h00}, /* 0xfbae */
            {8'h00}, /* 0xfbad */
            {8'h00}, /* 0xfbac */
            {8'h00}, /* 0xfbab */
            {8'h00}, /* 0xfbaa */
            {8'h00}, /* 0xfba9 */
            {8'h00}, /* 0xfba8 */
            {8'h00}, /* 0xfba7 */
            {8'h00}, /* 0xfba6 */
            {8'h00}, /* 0xfba5 */
            {8'h00}, /* 0xfba4 */
            {8'h00}, /* 0xfba3 */
            {8'h00}, /* 0xfba2 */
            {8'h00}, /* 0xfba1 */
            {8'h00}, /* 0xfba0 */
            {8'h00}, /* 0xfb9f */
            {8'h00}, /* 0xfb9e */
            {8'h00}, /* 0xfb9d */
            {8'h00}, /* 0xfb9c */
            {8'h00}, /* 0xfb9b */
            {8'h00}, /* 0xfb9a */
            {8'h00}, /* 0xfb99 */
            {8'h00}, /* 0xfb98 */
            {8'h00}, /* 0xfb97 */
            {8'h00}, /* 0xfb96 */
            {8'h00}, /* 0xfb95 */
            {8'h00}, /* 0xfb94 */
            {8'h00}, /* 0xfb93 */
            {8'h00}, /* 0xfb92 */
            {8'h00}, /* 0xfb91 */
            {8'h00}, /* 0xfb90 */
            {8'h00}, /* 0xfb8f */
            {8'h00}, /* 0xfb8e */
            {8'h00}, /* 0xfb8d */
            {8'h00}, /* 0xfb8c */
            {8'h00}, /* 0xfb8b */
            {8'h00}, /* 0xfb8a */
            {8'h00}, /* 0xfb89 */
            {8'h00}, /* 0xfb88 */
            {8'h00}, /* 0xfb87 */
            {8'h00}, /* 0xfb86 */
            {8'h00}, /* 0xfb85 */
            {8'h00}, /* 0xfb84 */
            {8'h00}, /* 0xfb83 */
            {8'h00}, /* 0xfb82 */
            {8'h00}, /* 0xfb81 */
            {8'h00}, /* 0xfb80 */
            {8'h00}, /* 0xfb7f */
            {8'h00}, /* 0xfb7e */
            {8'h00}, /* 0xfb7d */
            {8'h00}, /* 0xfb7c */
            {8'h00}, /* 0xfb7b */
            {8'h00}, /* 0xfb7a */
            {8'h00}, /* 0xfb79 */
            {8'h00}, /* 0xfb78 */
            {8'h00}, /* 0xfb77 */
            {8'h00}, /* 0xfb76 */
            {8'h00}, /* 0xfb75 */
            {8'h00}, /* 0xfb74 */
            {8'h00}, /* 0xfb73 */
            {8'h00}, /* 0xfb72 */
            {8'h00}, /* 0xfb71 */
            {8'h00}, /* 0xfb70 */
            {8'h00}, /* 0xfb6f */
            {8'h00}, /* 0xfb6e */
            {8'h00}, /* 0xfb6d */
            {8'h00}, /* 0xfb6c */
            {8'h00}, /* 0xfb6b */
            {8'h00}, /* 0xfb6a */
            {8'h00}, /* 0xfb69 */
            {8'h00}, /* 0xfb68 */
            {8'h00}, /* 0xfb67 */
            {8'h00}, /* 0xfb66 */
            {8'h00}, /* 0xfb65 */
            {8'h00}, /* 0xfb64 */
            {8'h00}, /* 0xfb63 */
            {8'h00}, /* 0xfb62 */
            {8'h00}, /* 0xfb61 */
            {8'h00}, /* 0xfb60 */
            {8'h00}, /* 0xfb5f */
            {8'h00}, /* 0xfb5e */
            {8'h00}, /* 0xfb5d */
            {8'h00}, /* 0xfb5c */
            {8'h00}, /* 0xfb5b */
            {8'h00}, /* 0xfb5a */
            {8'h00}, /* 0xfb59 */
            {8'h00}, /* 0xfb58 */
            {8'h00}, /* 0xfb57 */
            {8'h00}, /* 0xfb56 */
            {8'h00}, /* 0xfb55 */
            {8'h00}, /* 0xfb54 */
            {8'h00}, /* 0xfb53 */
            {8'h00}, /* 0xfb52 */
            {8'h00}, /* 0xfb51 */
            {8'h00}, /* 0xfb50 */
            {8'h00}, /* 0xfb4f */
            {8'h00}, /* 0xfb4e */
            {8'h00}, /* 0xfb4d */
            {8'h00}, /* 0xfb4c */
            {8'h00}, /* 0xfb4b */
            {8'h00}, /* 0xfb4a */
            {8'h00}, /* 0xfb49 */
            {8'h00}, /* 0xfb48 */
            {8'h00}, /* 0xfb47 */
            {8'h00}, /* 0xfb46 */
            {8'h00}, /* 0xfb45 */
            {8'h00}, /* 0xfb44 */
            {8'h00}, /* 0xfb43 */
            {8'h00}, /* 0xfb42 */
            {8'h00}, /* 0xfb41 */
            {8'h00}, /* 0xfb40 */
            {8'h00}, /* 0xfb3f */
            {8'h00}, /* 0xfb3e */
            {8'h00}, /* 0xfb3d */
            {8'h00}, /* 0xfb3c */
            {8'h00}, /* 0xfb3b */
            {8'h00}, /* 0xfb3a */
            {8'h00}, /* 0xfb39 */
            {8'h00}, /* 0xfb38 */
            {8'h00}, /* 0xfb37 */
            {8'h00}, /* 0xfb36 */
            {8'h00}, /* 0xfb35 */
            {8'h00}, /* 0xfb34 */
            {8'h00}, /* 0xfb33 */
            {8'h00}, /* 0xfb32 */
            {8'h00}, /* 0xfb31 */
            {8'h00}, /* 0xfb30 */
            {8'h00}, /* 0xfb2f */
            {8'h00}, /* 0xfb2e */
            {8'h00}, /* 0xfb2d */
            {8'h00}, /* 0xfb2c */
            {8'h00}, /* 0xfb2b */
            {8'h00}, /* 0xfb2a */
            {8'h00}, /* 0xfb29 */
            {8'h00}, /* 0xfb28 */
            {8'h00}, /* 0xfb27 */
            {8'h00}, /* 0xfb26 */
            {8'h00}, /* 0xfb25 */
            {8'h00}, /* 0xfb24 */
            {8'h00}, /* 0xfb23 */
            {8'h00}, /* 0xfb22 */
            {8'h00}, /* 0xfb21 */
            {8'h00}, /* 0xfb20 */
            {8'h00}, /* 0xfb1f */
            {8'h00}, /* 0xfb1e */
            {8'h00}, /* 0xfb1d */
            {8'h00}, /* 0xfb1c */
            {8'h00}, /* 0xfb1b */
            {8'h00}, /* 0xfb1a */
            {8'h00}, /* 0xfb19 */
            {8'h00}, /* 0xfb18 */
            {8'h00}, /* 0xfb17 */
            {8'h00}, /* 0xfb16 */
            {8'h00}, /* 0xfb15 */
            {8'h00}, /* 0xfb14 */
            {8'h00}, /* 0xfb13 */
            {8'h00}, /* 0xfb12 */
            {8'h00}, /* 0xfb11 */
            {8'h00}, /* 0xfb10 */
            {8'h00}, /* 0xfb0f */
            {8'h00}, /* 0xfb0e */
            {8'h00}, /* 0xfb0d */
            {8'h00}, /* 0xfb0c */
            {8'h00}, /* 0xfb0b */
            {8'h00}, /* 0xfb0a */
            {8'h00}, /* 0xfb09 */
            {8'h00}, /* 0xfb08 */
            {8'h00}, /* 0xfb07 */
            {8'h00}, /* 0xfb06 */
            {8'h00}, /* 0xfb05 */
            {8'h00}, /* 0xfb04 */
            {8'h00}, /* 0xfb03 */
            {8'h00}, /* 0xfb02 */
            {8'h00}, /* 0xfb01 */
            {8'h00}, /* 0xfb00 */
            {8'h00}, /* 0xfaff */
            {8'h00}, /* 0xfafe */
            {8'h00}, /* 0xfafd */
            {8'h00}, /* 0xfafc */
            {8'h00}, /* 0xfafb */
            {8'h00}, /* 0xfafa */
            {8'h00}, /* 0xfaf9 */
            {8'h00}, /* 0xfaf8 */
            {8'h00}, /* 0xfaf7 */
            {8'h00}, /* 0xfaf6 */
            {8'h00}, /* 0xfaf5 */
            {8'h00}, /* 0xfaf4 */
            {8'h00}, /* 0xfaf3 */
            {8'h00}, /* 0xfaf2 */
            {8'h00}, /* 0xfaf1 */
            {8'h00}, /* 0xfaf0 */
            {8'h00}, /* 0xfaef */
            {8'h00}, /* 0xfaee */
            {8'h00}, /* 0xfaed */
            {8'h00}, /* 0xfaec */
            {8'h00}, /* 0xfaeb */
            {8'h00}, /* 0xfaea */
            {8'h00}, /* 0xfae9 */
            {8'h00}, /* 0xfae8 */
            {8'h00}, /* 0xfae7 */
            {8'h00}, /* 0xfae6 */
            {8'h00}, /* 0xfae5 */
            {8'h00}, /* 0xfae4 */
            {8'h00}, /* 0xfae3 */
            {8'h00}, /* 0xfae2 */
            {8'h00}, /* 0xfae1 */
            {8'h00}, /* 0xfae0 */
            {8'h00}, /* 0xfadf */
            {8'h00}, /* 0xfade */
            {8'h00}, /* 0xfadd */
            {8'h00}, /* 0xfadc */
            {8'h00}, /* 0xfadb */
            {8'h00}, /* 0xfada */
            {8'h00}, /* 0xfad9 */
            {8'h00}, /* 0xfad8 */
            {8'h00}, /* 0xfad7 */
            {8'h00}, /* 0xfad6 */
            {8'h00}, /* 0xfad5 */
            {8'h00}, /* 0xfad4 */
            {8'h00}, /* 0xfad3 */
            {8'h00}, /* 0xfad2 */
            {8'h00}, /* 0xfad1 */
            {8'h00}, /* 0xfad0 */
            {8'h00}, /* 0xfacf */
            {8'h00}, /* 0xface */
            {8'h00}, /* 0xfacd */
            {8'h00}, /* 0xfacc */
            {8'h00}, /* 0xfacb */
            {8'h00}, /* 0xfaca */
            {8'h00}, /* 0xfac9 */
            {8'h00}, /* 0xfac8 */
            {8'h00}, /* 0xfac7 */
            {8'h00}, /* 0xfac6 */
            {8'h00}, /* 0xfac5 */
            {8'h00}, /* 0xfac4 */
            {8'h00}, /* 0xfac3 */
            {8'h00}, /* 0xfac2 */
            {8'h00}, /* 0xfac1 */
            {8'h00}, /* 0xfac0 */
            {8'h00}, /* 0xfabf */
            {8'h00}, /* 0xfabe */
            {8'h00}, /* 0xfabd */
            {8'h00}, /* 0xfabc */
            {8'h00}, /* 0xfabb */
            {8'h00}, /* 0xfaba */
            {8'h00}, /* 0xfab9 */
            {8'h00}, /* 0xfab8 */
            {8'h00}, /* 0xfab7 */
            {8'h00}, /* 0xfab6 */
            {8'h00}, /* 0xfab5 */
            {8'h00}, /* 0xfab4 */
            {8'h00}, /* 0xfab3 */
            {8'h00}, /* 0xfab2 */
            {8'h00}, /* 0xfab1 */
            {8'h00}, /* 0xfab0 */
            {8'h00}, /* 0xfaaf */
            {8'h00}, /* 0xfaae */
            {8'h00}, /* 0xfaad */
            {8'h00}, /* 0xfaac */
            {8'h00}, /* 0xfaab */
            {8'h00}, /* 0xfaaa */
            {8'h00}, /* 0xfaa9 */
            {8'h00}, /* 0xfaa8 */
            {8'h00}, /* 0xfaa7 */
            {8'h00}, /* 0xfaa6 */
            {8'h00}, /* 0xfaa5 */
            {8'h00}, /* 0xfaa4 */
            {8'h00}, /* 0xfaa3 */
            {8'h00}, /* 0xfaa2 */
            {8'h00}, /* 0xfaa1 */
            {8'h00}, /* 0xfaa0 */
            {8'h00}, /* 0xfa9f */
            {8'h00}, /* 0xfa9e */
            {8'h00}, /* 0xfa9d */
            {8'h00}, /* 0xfa9c */
            {8'h00}, /* 0xfa9b */
            {8'h00}, /* 0xfa9a */
            {8'h00}, /* 0xfa99 */
            {8'h00}, /* 0xfa98 */
            {8'h00}, /* 0xfa97 */
            {8'h00}, /* 0xfa96 */
            {8'h00}, /* 0xfa95 */
            {8'h00}, /* 0xfa94 */
            {8'h00}, /* 0xfa93 */
            {8'h00}, /* 0xfa92 */
            {8'h00}, /* 0xfa91 */
            {8'h00}, /* 0xfa90 */
            {8'h00}, /* 0xfa8f */
            {8'h00}, /* 0xfa8e */
            {8'h00}, /* 0xfa8d */
            {8'h00}, /* 0xfa8c */
            {8'h00}, /* 0xfa8b */
            {8'h00}, /* 0xfa8a */
            {8'h00}, /* 0xfa89 */
            {8'h00}, /* 0xfa88 */
            {8'h00}, /* 0xfa87 */
            {8'h00}, /* 0xfa86 */
            {8'h00}, /* 0xfa85 */
            {8'h00}, /* 0xfa84 */
            {8'h00}, /* 0xfa83 */
            {8'h00}, /* 0xfa82 */
            {8'h00}, /* 0xfa81 */
            {8'h00}, /* 0xfa80 */
            {8'h00}, /* 0xfa7f */
            {8'h00}, /* 0xfa7e */
            {8'h00}, /* 0xfa7d */
            {8'h00}, /* 0xfa7c */
            {8'h00}, /* 0xfa7b */
            {8'h00}, /* 0xfa7a */
            {8'h00}, /* 0xfa79 */
            {8'h00}, /* 0xfa78 */
            {8'h00}, /* 0xfa77 */
            {8'h00}, /* 0xfa76 */
            {8'h00}, /* 0xfa75 */
            {8'h00}, /* 0xfa74 */
            {8'h00}, /* 0xfa73 */
            {8'h00}, /* 0xfa72 */
            {8'h00}, /* 0xfa71 */
            {8'h00}, /* 0xfa70 */
            {8'h00}, /* 0xfa6f */
            {8'h00}, /* 0xfa6e */
            {8'h00}, /* 0xfa6d */
            {8'h00}, /* 0xfa6c */
            {8'h00}, /* 0xfa6b */
            {8'h00}, /* 0xfa6a */
            {8'h00}, /* 0xfa69 */
            {8'h00}, /* 0xfa68 */
            {8'h00}, /* 0xfa67 */
            {8'h00}, /* 0xfa66 */
            {8'h00}, /* 0xfa65 */
            {8'h00}, /* 0xfa64 */
            {8'h00}, /* 0xfa63 */
            {8'h00}, /* 0xfa62 */
            {8'h00}, /* 0xfa61 */
            {8'h00}, /* 0xfa60 */
            {8'h00}, /* 0xfa5f */
            {8'h00}, /* 0xfa5e */
            {8'h00}, /* 0xfa5d */
            {8'h00}, /* 0xfa5c */
            {8'h00}, /* 0xfa5b */
            {8'h00}, /* 0xfa5a */
            {8'h00}, /* 0xfa59 */
            {8'h00}, /* 0xfa58 */
            {8'h00}, /* 0xfa57 */
            {8'h00}, /* 0xfa56 */
            {8'h00}, /* 0xfa55 */
            {8'h00}, /* 0xfa54 */
            {8'h00}, /* 0xfa53 */
            {8'h00}, /* 0xfa52 */
            {8'h00}, /* 0xfa51 */
            {8'h00}, /* 0xfa50 */
            {8'h00}, /* 0xfa4f */
            {8'h00}, /* 0xfa4e */
            {8'h00}, /* 0xfa4d */
            {8'h00}, /* 0xfa4c */
            {8'h00}, /* 0xfa4b */
            {8'h00}, /* 0xfa4a */
            {8'h00}, /* 0xfa49 */
            {8'h00}, /* 0xfa48 */
            {8'h00}, /* 0xfa47 */
            {8'h00}, /* 0xfa46 */
            {8'h00}, /* 0xfa45 */
            {8'h00}, /* 0xfa44 */
            {8'h00}, /* 0xfa43 */
            {8'h00}, /* 0xfa42 */
            {8'h00}, /* 0xfa41 */
            {8'h00}, /* 0xfa40 */
            {8'h00}, /* 0xfa3f */
            {8'h00}, /* 0xfa3e */
            {8'h00}, /* 0xfa3d */
            {8'h00}, /* 0xfa3c */
            {8'h00}, /* 0xfa3b */
            {8'h00}, /* 0xfa3a */
            {8'h00}, /* 0xfa39 */
            {8'h00}, /* 0xfa38 */
            {8'h00}, /* 0xfa37 */
            {8'h00}, /* 0xfa36 */
            {8'h00}, /* 0xfa35 */
            {8'h00}, /* 0xfa34 */
            {8'h00}, /* 0xfa33 */
            {8'h00}, /* 0xfa32 */
            {8'h00}, /* 0xfa31 */
            {8'h00}, /* 0xfa30 */
            {8'h00}, /* 0xfa2f */
            {8'h00}, /* 0xfa2e */
            {8'h00}, /* 0xfa2d */
            {8'h00}, /* 0xfa2c */
            {8'h00}, /* 0xfa2b */
            {8'h00}, /* 0xfa2a */
            {8'h00}, /* 0xfa29 */
            {8'h00}, /* 0xfa28 */
            {8'h00}, /* 0xfa27 */
            {8'h00}, /* 0xfa26 */
            {8'h00}, /* 0xfa25 */
            {8'h00}, /* 0xfa24 */
            {8'h00}, /* 0xfa23 */
            {8'h00}, /* 0xfa22 */
            {8'h00}, /* 0xfa21 */
            {8'h00}, /* 0xfa20 */
            {8'h00}, /* 0xfa1f */
            {8'h00}, /* 0xfa1e */
            {8'h00}, /* 0xfa1d */
            {8'h00}, /* 0xfa1c */
            {8'h00}, /* 0xfa1b */
            {8'h00}, /* 0xfa1a */
            {8'h00}, /* 0xfa19 */
            {8'h00}, /* 0xfa18 */
            {8'h00}, /* 0xfa17 */
            {8'h00}, /* 0xfa16 */
            {8'h00}, /* 0xfa15 */
            {8'h00}, /* 0xfa14 */
            {8'h00}, /* 0xfa13 */
            {8'h00}, /* 0xfa12 */
            {8'h00}, /* 0xfa11 */
            {8'h00}, /* 0xfa10 */
            {8'h00}, /* 0xfa0f */
            {8'h00}, /* 0xfa0e */
            {8'h00}, /* 0xfa0d */
            {8'h00}, /* 0xfa0c */
            {8'h00}, /* 0xfa0b */
            {8'h00}, /* 0xfa0a */
            {8'h00}, /* 0xfa09 */
            {8'h00}, /* 0xfa08 */
            {8'h00}, /* 0xfa07 */
            {8'h00}, /* 0xfa06 */
            {8'h00}, /* 0xfa05 */
            {8'h00}, /* 0xfa04 */
            {8'h00}, /* 0xfa03 */
            {8'h00}, /* 0xfa02 */
            {8'h00}, /* 0xfa01 */
            {8'h00}, /* 0xfa00 */
            {8'h00}, /* 0xf9ff */
            {8'h00}, /* 0xf9fe */
            {8'h00}, /* 0xf9fd */
            {8'h00}, /* 0xf9fc */
            {8'h00}, /* 0xf9fb */
            {8'h00}, /* 0xf9fa */
            {8'h00}, /* 0xf9f9 */
            {8'h00}, /* 0xf9f8 */
            {8'h00}, /* 0xf9f7 */
            {8'h00}, /* 0xf9f6 */
            {8'h00}, /* 0xf9f5 */
            {8'h00}, /* 0xf9f4 */
            {8'h00}, /* 0xf9f3 */
            {8'h00}, /* 0xf9f2 */
            {8'h00}, /* 0xf9f1 */
            {8'h00}, /* 0xf9f0 */
            {8'h00}, /* 0xf9ef */
            {8'h00}, /* 0xf9ee */
            {8'h00}, /* 0xf9ed */
            {8'h00}, /* 0xf9ec */
            {8'h00}, /* 0xf9eb */
            {8'h00}, /* 0xf9ea */
            {8'h00}, /* 0xf9e9 */
            {8'h00}, /* 0xf9e8 */
            {8'h00}, /* 0xf9e7 */
            {8'h00}, /* 0xf9e6 */
            {8'h00}, /* 0xf9e5 */
            {8'h00}, /* 0xf9e4 */
            {8'h00}, /* 0xf9e3 */
            {8'h00}, /* 0xf9e2 */
            {8'h00}, /* 0xf9e1 */
            {8'h00}, /* 0xf9e0 */
            {8'h00}, /* 0xf9df */
            {8'h00}, /* 0xf9de */
            {8'h00}, /* 0xf9dd */
            {8'h00}, /* 0xf9dc */
            {8'h00}, /* 0xf9db */
            {8'h00}, /* 0xf9da */
            {8'h00}, /* 0xf9d9 */
            {8'h00}, /* 0xf9d8 */
            {8'h00}, /* 0xf9d7 */
            {8'h00}, /* 0xf9d6 */
            {8'h00}, /* 0xf9d5 */
            {8'h00}, /* 0xf9d4 */
            {8'h00}, /* 0xf9d3 */
            {8'h00}, /* 0xf9d2 */
            {8'h00}, /* 0xf9d1 */
            {8'h00}, /* 0xf9d0 */
            {8'h00}, /* 0xf9cf */
            {8'h00}, /* 0xf9ce */
            {8'h00}, /* 0xf9cd */
            {8'h00}, /* 0xf9cc */
            {8'h00}, /* 0xf9cb */
            {8'h00}, /* 0xf9ca */
            {8'h00}, /* 0xf9c9 */
            {8'h00}, /* 0xf9c8 */
            {8'h00}, /* 0xf9c7 */
            {8'h00}, /* 0xf9c6 */
            {8'h00}, /* 0xf9c5 */
            {8'h00}, /* 0xf9c4 */
            {8'h00}, /* 0xf9c3 */
            {8'h00}, /* 0xf9c2 */
            {8'h00}, /* 0xf9c1 */
            {8'h00}, /* 0xf9c0 */
            {8'h00}, /* 0xf9bf */
            {8'h00}, /* 0xf9be */
            {8'h00}, /* 0xf9bd */
            {8'h00}, /* 0xf9bc */
            {8'h00}, /* 0xf9bb */
            {8'h00}, /* 0xf9ba */
            {8'h00}, /* 0xf9b9 */
            {8'h00}, /* 0xf9b8 */
            {8'h00}, /* 0xf9b7 */
            {8'h00}, /* 0xf9b6 */
            {8'h00}, /* 0xf9b5 */
            {8'h00}, /* 0xf9b4 */
            {8'h00}, /* 0xf9b3 */
            {8'h00}, /* 0xf9b2 */
            {8'h00}, /* 0xf9b1 */
            {8'h00}, /* 0xf9b0 */
            {8'h00}, /* 0xf9af */
            {8'h00}, /* 0xf9ae */
            {8'h00}, /* 0xf9ad */
            {8'h00}, /* 0xf9ac */
            {8'h00}, /* 0xf9ab */
            {8'h00}, /* 0xf9aa */
            {8'h00}, /* 0xf9a9 */
            {8'h00}, /* 0xf9a8 */
            {8'h00}, /* 0xf9a7 */
            {8'h00}, /* 0xf9a6 */
            {8'h00}, /* 0xf9a5 */
            {8'h00}, /* 0xf9a4 */
            {8'h00}, /* 0xf9a3 */
            {8'h00}, /* 0xf9a2 */
            {8'h00}, /* 0xf9a1 */
            {8'h00}, /* 0xf9a0 */
            {8'h00}, /* 0xf99f */
            {8'h00}, /* 0xf99e */
            {8'h00}, /* 0xf99d */
            {8'h00}, /* 0xf99c */
            {8'h00}, /* 0xf99b */
            {8'h00}, /* 0xf99a */
            {8'h00}, /* 0xf999 */
            {8'h00}, /* 0xf998 */
            {8'h00}, /* 0xf997 */
            {8'h00}, /* 0xf996 */
            {8'h00}, /* 0xf995 */
            {8'h00}, /* 0xf994 */
            {8'h00}, /* 0xf993 */
            {8'h00}, /* 0xf992 */
            {8'h00}, /* 0xf991 */
            {8'h00}, /* 0xf990 */
            {8'h00}, /* 0xf98f */
            {8'h00}, /* 0xf98e */
            {8'h00}, /* 0xf98d */
            {8'h00}, /* 0xf98c */
            {8'h00}, /* 0xf98b */
            {8'h00}, /* 0xf98a */
            {8'h00}, /* 0xf989 */
            {8'h00}, /* 0xf988 */
            {8'h00}, /* 0xf987 */
            {8'h00}, /* 0xf986 */
            {8'h00}, /* 0xf985 */
            {8'h00}, /* 0xf984 */
            {8'h00}, /* 0xf983 */
            {8'h00}, /* 0xf982 */
            {8'h00}, /* 0xf981 */
            {8'h00}, /* 0xf980 */
            {8'h00}, /* 0xf97f */
            {8'h00}, /* 0xf97e */
            {8'h00}, /* 0xf97d */
            {8'h00}, /* 0xf97c */
            {8'h00}, /* 0xf97b */
            {8'h00}, /* 0xf97a */
            {8'h00}, /* 0xf979 */
            {8'h00}, /* 0xf978 */
            {8'h00}, /* 0xf977 */
            {8'h00}, /* 0xf976 */
            {8'h00}, /* 0xf975 */
            {8'h00}, /* 0xf974 */
            {8'h00}, /* 0xf973 */
            {8'h00}, /* 0xf972 */
            {8'h00}, /* 0xf971 */
            {8'h00}, /* 0xf970 */
            {8'h00}, /* 0xf96f */
            {8'h00}, /* 0xf96e */
            {8'h00}, /* 0xf96d */
            {8'h00}, /* 0xf96c */
            {8'h00}, /* 0xf96b */
            {8'h00}, /* 0xf96a */
            {8'h00}, /* 0xf969 */
            {8'h00}, /* 0xf968 */
            {8'h00}, /* 0xf967 */
            {8'h00}, /* 0xf966 */
            {8'h00}, /* 0xf965 */
            {8'h00}, /* 0xf964 */
            {8'h00}, /* 0xf963 */
            {8'h00}, /* 0xf962 */
            {8'h00}, /* 0xf961 */
            {8'h00}, /* 0xf960 */
            {8'h00}, /* 0xf95f */
            {8'h00}, /* 0xf95e */
            {8'h00}, /* 0xf95d */
            {8'h00}, /* 0xf95c */
            {8'h00}, /* 0xf95b */
            {8'h00}, /* 0xf95a */
            {8'h00}, /* 0xf959 */
            {8'h00}, /* 0xf958 */
            {8'h00}, /* 0xf957 */
            {8'h00}, /* 0xf956 */
            {8'h00}, /* 0xf955 */
            {8'h00}, /* 0xf954 */
            {8'h00}, /* 0xf953 */
            {8'h00}, /* 0xf952 */
            {8'h00}, /* 0xf951 */
            {8'h00}, /* 0xf950 */
            {8'h00}, /* 0xf94f */
            {8'h00}, /* 0xf94e */
            {8'h00}, /* 0xf94d */
            {8'h00}, /* 0xf94c */
            {8'h00}, /* 0xf94b */
            {8'h00}, /* 0xf94a */
            {8'h00}, /* 0xf949 */
            {8'h00}, /* 0xf948 */
            {8'h00}, /* 0xf947 */
            {8'h00}, /* 0xf946 */
            {8'h00}, /* 0xf945 */
            {8'h00}, /* 0xf944 */
            {8'h00}, /* 0xf943 */
            {8'h00}, /* 0xf942 */
            {8'h00}, /* 0xf941 */
            {8'h00}, /* 0xf940 */
            {8'h00}, /* 0xf93f */
            {8'h00}, /* 0xf93e */
            {8'h00}, /* 0xf93d */
            {8'h00}, /* 0xf93c */
            {8'h00}, /* 0xf93b */
            {8'h00}, /* 0xf93a */
            {8'h00}, /* 0xf939 */
            {8'h00}, /* 0xf938 */
            {8'h00}, /* 0xf937 */
            {8'h00}, /* 0xf936 */
            {8'h00}, /* 0xf935 */
            {8'h00}, /* 0xf934 */
            {8'h00}, /* 0xf933 */
            {8'h00}, /* 0xf932 */
            {8'h00}, /* 0xf931 */
            {8'h00}, /* 0xf930 */
            {8'h00}, /* 0xf92f */
            {8'h00}, /* 0xf92e */
            {8'h00}, /* 0xf92d */
            {8'h00}, /* 0xf92c */
            {8'h00}, /* 0xf92b */
            {8'h00}, /* 0xf92a */
            {8'h00}, /* 0xf929 */
            {8'h00}, /* 0xf928 */
            {8'h00}, /* 0xf927 */
            {8'h00}, /* 0xf926 */
            {8'h00}, /* 0xf925 */
            {8'h00}, /* 0xf924 */
            {8'h00}, /* 0xf923 */
            {8'h00}, /* 0xf922 */
            {8'h00}, /* 0xf921 */
            {8'h00}, /* 0xf920 */
            {8'h00}, /* 0xf91f */
            {8'h00}, /* 0xf91e */
            {8'h00}, /* 0xf91d */
            {8'h00}, /* 0xf91c */
            {8'h00}, /* 0xf91b */
            {8'h00}, /* 0xf91a */
            {8'h00}, /* 0xf919 */
            {8'h00}, /* 0xf918 */
            {8'h00}, /* 0xf917 */
            {8'h00}, /* 0xf916 */
            {8'h00}, /* 0xf915 */
            {8'h00}, /* 0xf914 */
            {8'h00}, /* 0xf913 */
            {8'h00}, /* 0xf912 */
            {8'h00}, /* 0xf911 */
            {8'h00}, /* 0xf910 */
            {8'h00}, /* 0xf90f */
            {8'h00}, /* 0xf90e */
            {8'h00}, /* 0xf90d */
            {8'h00}, /* 0xf90c */
            {8'h00}, /* 0xf90b */
            {8'h00}, /* 0xf90a */
            {8'h00}, /* 0xf909 */
            {8'h00}, /* 0xf908 */
            {8'h00}, /* 0xf907 */
            {8'h00}, /* 0xf906 */
            {8'h00}, /* 0xf905 */
            {8'h00}, /* 0xf904 */
            {8'h00}, /* 0xf903 */
            {8'h00}, /* 0xf902 */
            {8'h00}, /* 0xf901 */
            {8'h00}, /* 0xf900 */
            {8'h00}, /* 0xf8ff */
            {8'h00}, /* 0xf8fe */
            {8'h00}, /* 0xf8fd */
            {8'h00}, /* 0xf8fc */
            {8'h00}, /* 0xf8fb */
            {8'h00}, /* 0xf8fa */
            {8'h00}, /* 0xf8f9 */
            {8'h00}, /* 0xf8f8 */
            {8'h00}, /* 0xf8f7 */
            {8'h00}, /* 0xf8f6 */
            {8'h00}, /* 0xf8f5 */
            {8'h00}, /* 0xf8f4 */
            {8'h00}, /* 0xf8f3 */
            {8'h00}, /* 0xf8f2 */
            {8'h00}, /* 0xf8f1 */
            {8'h00}, /* 0xf8f0 */
            {8'h00}, /* 0xf8ef */
            {8'h00}, /* 0xf8ee */
            {8'h00}, /* 0xf8ed */
            {8'h00}, /* 0xf8ec */
            {8'h00}, /* 0xf8eb */
            {8'h00}, /* 0xf8ea */
            {8'h00}, /* 0xf8e9 */
            {8'h00}, /* 0xf8e8 */
            {8'h00}, /* 0xf8e7 */
            {8'h00}, /* 0xf8e6 */
            {8'h00}, /* 0xf8e5 */
            {8'h00}, /* 0xf8e4 */
            {8'h00}, /* 0xf8e3 */
            {8'h00}, /* 0xf8e2 */
            {8'h00}, /* 0xf8e1 */
            {8'h00}, /* 0xf8e0 */
            {8'h00}, /* 0xf8df */
            {8'h00}, /* 0xf8de */
            {8'h00}, /* 0xf8dd */
            {8'h00}, /* 0xf8dc */
            {8'h00}, /* 0xf8db */
            {8'h00}, /* 0xf8da */
            {8'h00}, /* 0xf8d9 */
            {8'h00}, /* 0xf8d8 */
            {8'h00}, /* 0xf8d7 */
            {8'h00}, /* 0xf8d6 */
            {8'h00}, /* 0xf8d5 */
            {8'h00}, /* 0xf8d4 */
            {8'h00}, /* 0xf8d3 */
            {8'h00}, /* 0xf8d2 */
            {8'h00}, /* 0xf8d1 */
            {8'h00}, /* 0xf8d0 */
            {8'h00}, /* 0xf8cf */
            {8'h00}, /* 0xf8ce */
            {8'h00}, /* 0xf8cd */
            {8'h00}, /* 0xf8cc */
            {8'h00}, /* 0xf8cb */
            {8'h00}, /* 0xf8ca */
            {8'h00}, /* 0xf8c9 */
            {8'h00}, /* 0xf8c8 */
            {8'h00}, /* 0xf8c7 */
            {8'h00}, /* 0xf8c6 */
            {8'h00}, /* 0xf8c5 */
            {8'h00}, /* 0xf8c4 */
            {8'h00}, /* 0xf8c3 */
            {8'h00}, /* 0xf8c2 */
            {8'h00}, /* 0xf8c1 */
            {8'h00}, /* 0xf8c0 */
            {8'h00}, /* 0xf8bf */
            {8'h00}, /* 0xf8be */
            {8'h00}, /* 0xf8bd */
            {8'h00}, /* 0xf8bc */
            {8'h00}, /* 0xf8bb */
            {8'h00}, /* 0xf8ba */
            {8'h00}, /* 0xf8b9 */
            {8'h00}, /* 0xf8b8 */
            {8'h00}, /* 0xf8b7 */
            {8'h00}, /* 0xf8b6 */
            {8'h00}, /* 0xf8b5 */
            {8'h00}, /* 0xf8b4 */
            {8'h00}, /* 0xf8b3 */
            {8'h00}, /* 0xf8b2 */
            {8'h00}, /* 0xf8b1 */
            {8'h00}, /* 0xf8b0 */
            {8'h00}, /* 0xf8af */
            {8'h00}, /* 0xf8ae */
            {8'h00}, /* 0xf8ad */
            {8'h00}, /* 0xf8ac */
            {8'h00}, /* 0xf8ab */
            {8'h00}, /* 0xf8aa */
            {8'h00}, /* 0xf8a9 */
            {8'h00}, /* 0xf8a8 */
            {8'h00}, /* 0xf8a7 */
            {8'h00}, /* 0xf8a6 */
            {8'h00}, /* 0xf8a5 */
            {8'h00}, /* 0xf8a4 */
            {8'h00}, /* 0xf8a3 */
            {8'h00}, /* 0xf8a2 */
            {8'h00}, /* 0xf8a1 */
            {8'h00}, /* 0xf8a0 */
            {8'h00}, /* 0xf89f */
            {8'h00}, /* 0xf89e */
            {8'h00}, /* 0xf89d */
            {8'h00}, /* 0xf89c */
            {8'h00}, /* 0xf89b */
            {8'h00}, /* 0xf89a */
            {8'h00}, /* 0xf899 */
            {8'h00}, /* 0xf898 */
            {8'h00}, /* 0xf897 */
            {8'h00}, /* 0xf896 */
            {8'h00}, /* 0xf895 */
            {8'h00}, /* 0xf894 */
            {8'h00}, /* 0xf893 */
            {8'h00}, /* 0xf892 */
            {8'h00}, /* 0xf891 */
            {8'h00}, /* 0xf890 */
            {8'h00}, /* 0xf88f */
            {8'h00}, /* 0xf88e */
            {8'h00}, /* 0xf88d */
            {8'h00}, /* 0xf88c */
            {8'h00}, /* 0xf88b */
            {8'h00}, /* 0xf88a */
            {8'h00}, /* 0xf889 */
            {8'h00}, /* 0xf888 */
            {8'h00}, /* 0xf887 */
            {8'h00}, /* 0xf886 */
            {8'h00}, /* 0xf885 */
            {8'h00}, /* 0xf884 */
            {8'h00}, /* 0xf883 */
            {8'h00}, /* 0xf882 */
            {8'h00}, /* 0xf881 */
            {8'h00}, /* 0xf880 */
            {8'h00}, /* 0xf87f */
            {8'h00}, /* 0xf87e */
            {8'h00}, /* 0xf87d */
            {8'h00}, /* 0xf87c */
            {8'h00}, /* 0xf87b */
            {8'h00}, /* 0xf87a */
            {8'h00}, /* 0xf879 */
            {8'h00}, /* 0xf878 */
            {8'h00}, /* 0xf877 */
            {8'h00}, /* 0xf876 */
            {8'h00}, /* 0xf875 */
            {8'h00}, /* 0xf874 */
            {8'h00}, /* 0xf873 */
            {8'h00}, /* 0xf872 */
            {8'h00}, /* 0xf871 */
            {8'h00}, /* 0xf870 */
            {8'h00}, /* 0xf86f */
            {8'h00}, /* 0xf86e */
            {8'h00}, /* 0xf86d */
            {8'h00}, /* 0xf86c */
            {8'h00}, /* 0xf86b */
            {8'h00}, /* 0xf86a */
            {8'h00}, /* 0xf869 */
            {8'h00}, /* 0xf868 */
            {8'h00}, /* 0xf867 */
            {8'h00}, /* 0xf866 */
            {8'h00}, /* 0xf865 */
            {8'h00}, /* 0xf864 */
            {8'h00}, /* 0xf863 */
            {8'h00}, /* 0xf862 */
            {8'h00}, /* 0xf861 */
            {8'h00}, /* 0xf860 */
            {8'h00}, /* 0xf85f */
            {8'h00}, /* 0xf85e */
            {8'h00}, /* 0xf85d */
            {8'h00}, /* 0xf85c */
            {8'h00}, /* 0xf85b */
            {8'h00}, /* 0xf85a */
            {8'h00}, /* 0xf859 */
            {8'h00}, /* 0xf858 */
            {8'h00}, /* 0xf857 */
            {8'h00}, /* 0xf856 */
            {8'h00}, /* 0xf855 */
            {8'h00}, /* 0xf854 */
            {8'h00}, /* 0xf853 */
            {8'h00}, /* 0xf852 */
            {8'h00}, /* 0xf851 */
            {8'h00}, /* 0xf850 */
            {8'h00}, /* 0xf84f */
            {8'h00}, /* 0xf84e */
            {8'h00}, /* 0xf84d */
            {8'h00}, /* 0xf84c */
            {8'h00}, /* 0xf84b */
            {8'h00}, /* 0xf84a */
            {8'h00}, /* 0xf849 */
            {8'h00}, /* 0xf848 */
            {8'h00}, /* 0xf847 */
            {8'h00}, /* 0xf846 */
            {8'h00}, /* 0xf845 */
            {8'h00}, /* 0xf844 */
            {8'h00}, /* 0xf843 */
            {8'h00}, /* 0xf842 */
            {8'h00}, /* 0xf841 */
            {8'h00}, /* 0xf840 */
            {8'h00}, /* 0xf83f */
            {8'h00}, /* 0xf83e */
            {8'h00}, /* 0xf83d */
            {8'h00}, /* 0xf83c */
            {8'h00}, /* 0xf83b */
            {8'h00}, /* 0xf83a */
            {8'h00}, /* 0xf839 */
            {8'h00}, /* 0xf838 */
            {8'h00}, /* 0xf837 */
            {8'h00}, /* 0xf836 */
            {8'h00}, /* 0xf835 */
            {8'h00}, /* 0xf834 */
            {8'h00}, /* 0xf833 */
            {8'h00}, /* 0xf832 */
            {8'h00}, /* 0xf831 */
            {8'h00}, /* 0xf830 */
            {8'h00}, /* 0xf82f */
            {8'h00}, /* 0xf82e */
            {8'h00}, /* 0xf82d */
            {8'h00}, /* 0xf82c */
            {8'h00}, /* 0xf82b */
            {8'h00}, /* 0xf82a */
            {8'h00}, /* 0xf829 */
            {8'h00}, /* 0xf828 */
            {8'h00}, /* 0xf827 */
            {8'h00}, /* 0xf826 */
            {8'h00}, /* 0xf825 */
            {8'h00}, /* 0xf824 */
            {8'h00}, /* 0xf823 */
            {8'h00}, /* 0xf822 */
            {8'h00}, /* 0xf821 */
            {8'h00}, /* 0xf820 */
            {8'h00}, /* 0xf81f */
            {8'h00}, /* 0xf81e */
            {8'h00}, /* 0xf81d */
            {8'h00}, /* 0xf81c */
            {8'h00}, /* 0xf81b */
            {8'h00}, /* 0xf81a */
            {8'h00}, /* 0xf819 */
            {8'h00}, /* 0xf818 */
            {8'h00}, /* 0xf817 */
            {8'h00}, /* 0xf816 */
            {8'h00}, /* 0xf815 */
            {8'h00}, /* 0xf814 */
            {8'h00}, /* 0xf813 */
            {8'h00}, /* 0xf812 */
            {8'h00}, /* 0xf811 */
            {8'h00}, /* 0xf810 */
            {8'h00}, /* 0xf80f */
            {8'h00}, /* 0xf80e */
            {8'h00}, /* 0xf80d */
            {8'h00}, /* 0xf80c */
            {8'h00}, /* 0xf80b */
            {8'h00}, /* 0xf80a */
            {8'h00}, /* 0xf809 */
            {8'h00}, /* 0xf808 */
            {8'h00}, /* 0xf807 */
            {8'h00}, /* 0xf806 */
            {8'h00}, /* 0xf805 */
            {8'h00}, /* 0xf804 */
            {8'h00}, /* 0xf803 */
            {8'h00}, /* 0xf802 */
            {8'h00}, /* 0xf801 */
            {8'h00}, /* 0xf800 */
            {8'h00}, /* 0xf7ff */
            {8'h00}, /* 0xf7fe */
            {8'h00}, /* 0xf7fd */
            {8'h00}, /* 0xf7fc */
            {8'h00}, /* 0xf7fb */
            {8'h00}, /* 0xf7fa */
            {8'h00}, /* 0xf7f9 */
            {8'h00}, /* 0xf7f8 */
            {8'h00}, /* 0xf7f7 */
            {8'h00}, /* 0xf7f6 */
            {8'h00}, /* 0xf7f5 */
            {8'h00}, /* 0xf7f4 */
            {8'h00}, /* 0xf7f3 */
            {8'h00}, /* 0xf7f2 */
            {8'h00}, /* 0xf7f1 */
            {8'h00}, /* 0xf7f0 */
            {8'h00}, /* 0xf7ef */
            {8'h00}, /* 0xf7ee */
            {8'h00}, /* 0xf7ed */
            {8'h00}, /* 0xf7ec */
            {8'h00}, /* 0xf7eb */
            {8'h00}, /* 0xf7ea */
            {8'h00}, /* 0xf7e9 */
            {8'h00}, /* 0xf7e8 */
            {8'h00}, /* 0xf7e7 */
            {8'h00}, /* 0xf7e6 */
            {8'h00}, /* 0xf7e5 */
            {8'h00}, /* 0xf7e4 */
            {8'h00}, /* 0xf7e3 */
            {8'h00}, /* 0xf7e2 */
            {8'h00}, /* 0xf7e1 */
            {8'h00}, /* 0xf7e0 */
            {8'h00}, /* 0xf7df */
            {8'h00}, /* 0xf7de */
            {8'h00}, /* 0xf7dd */
            {8'h00}, /* 0xf7dc */
            {8'h00}, /* 0xf7db */
            {8'h00}, /* 0xf7da */
            {8'h00}, /* 0xf7d9 */
            {8'h00}, /* 0xf7d8 */
            {8'h00}, /* 0xf7d7 */
            {8'h00}, /* 0xf7d6 */
            {8'h00}, /* 0xf7d5 */
            {8'h00}, /* 0xf7d4 */
            {8'h00}, /* 0xf7d3 */
            {8'h00}, /* 0xf7d2 */
            {8'h00}, /* 0xf7d1 */
            {8'h00}, /* 0xf7d0 */
            {8'h00}, /* 0xf7cf */
            {8'h00}, /* 0xf7ce */
            {8'h00}, /* 0xf7cd */
            {8'h00}, /* 0xf7cc */
            {8'h00}, /* 0xf7cb */
            {8'h00}, /* 0xf7ca */
            {8'h00}, /* 0xf7c9 */
            {8'h00}, /* 0xf7c8 */
            {8'h00}, /* 0xf7c7 */
            {8'h00}, /* 0xf7c6 */
            {8'h00}, /* 0xf7c5 */
            {8'h00}, /* 0xf7c4 */
            {8'h00}, /* 0xf7c3 */
            {8'h00}, /* 0xf7c2 */
            {8'h00}, /* 0xf7c1 */
            {8'h00}, /* 0xf7c0 */
            {8'h00}, /* 0xf7bf */
            {8'h00}, /* 0xf7be */
            {8'h00}, /* 0xf7bd */
            {8'h00}, /* 0xf7bc */
            {8'h00}, /* 0xf7bb */
            {8'h00}, /* 0xf7ba */
            {8'h00}, /* 0xf7b9 */
            {8'h00}, /* 0xf7b8 */
            {8'h00}, /* 0xf7b7 */
            {8'h00}, /* 0xf7b6 */
            {8'h00}, /* 0xf7b5 */
            {8'h00}, /* 0xf7b4 */
            {8'h00}, /* 0xf7b3 */
            {8'h00}, /* 0xf7b2 */
            {8'h00}, /* 0xf7b1 */
            {8'h00}, /* 0xf7b0 */
            {8'h00}, /* 0xf7af */
            {8'h00}, /* 0xf7ae */
            {8'h00}, /* 0xf7ad */
            {8'h00}, /* 0xf7ac */
            {8'h00}, /* 0xf7ab */
            {8'h00}, /* 0xf7aa */
            {8'h00}, /* 0xf7a9 */
            {8'h00}, /* 0xf7a8 */
            {8'h00}, /* 0xf7a7 */
            {8'h00}, /* 0xf7a6 */
            {8'h00}, /* 0xf7a5 */
            {8'h00}, /* 0xf7a4 */
            {8'h00}, /* 0xf7a3 */
            {8'h00}, /* 0xf7a2 */
            {8'h00}, /* 0xf7a1 */
            {8'h00}, /* 0xf7a0 */
            {8'h00}, /* 0xf79f */
            {8'h00}, /* 0xf79e */
            {8'h00}, /* 0xf79d */
            {8'h00}, /* 0xf79c */
            {8'h00}, /* 0xf79b */
            {8'h00}, /* 0xf79a */
            {8'h00}, /* 0xf799 */
            {8'h00}, /* 0xf798 */
            {8'h00}, /* 0xf797 */
            {8'h00}, /* 0xf796 */
            {8'h00}, /* 0xf795 */
            {8'h00}, /* 0xf794 */
            {8'h00}, /* 0xf793 */
            {8'h00}, /* 0xf792 */
            {8'h00}, /* 0xf791 */
            {8'h00}, /* 0xf790 */
            {8'h00}, /* 0xf78f */
            {8'h00}, /* 0xf78e */
            {8'h00}, /* 0xf78d */
            {8'h00}, /* 0xf78c */
            {8'h00}, /* 0xf78b */
            {8'h00}, /* 0xf78a */
            {8'h00}, /* 0xf789 */
            {8'h00}, /* 0xf788 */
            {8'h00}, /* 0xf787 */
            {8'h00}, /* 0xf786 */
            {8'h00}, /* 0xf785 */
            {8'h00}, /* 0xf784 */
            {8'h00}, /* 0xf783 */
            {8'h00}, /* 0xf782 */
            {8'h00}, /* 0xf781 */
            {8'h00}, /* 0xf780 */
            {8'h00}, /* 0xf77f */
            {8'h00}, /* 0xf77e */
            {8'h00}, /* 0xf77d */
            {8'h00}, /* 0xf77c */
            {8'h00}, /* 0xf77b */
            {8'h00}, /* 0xf77a */
            {8'h00}, /* 0xf779 */
            {8'h00}, /* 0xf778 */
            {8'h00}, /* 0xf777 */
            {8'h00}, /* 0xf776 */
            {8'h00}, /* 0xf775 */
            {8'h00}, /* 0xf774 */
            {8'h00}, /* 0xf773 */
            {8'h00}, /* 0xf772 */
            {8'h00}, /* 0xf771 */
            {8'h00}, /* 0xf770 */
            {8'h00}, /* 0xf76f */
            {8'h00}, /* 0xf76e */
            {8'h00}, /* 0xf76d */
            {8'h00}, /* 0xf76c */
            {8'h00}, /* 0xf76b */
            {8'h00}, /* 0xf76a */
            {8'h00}, /* 0xf769 */
            {8'h00}, /* 0xf768 */
            {8'h00}, /* 0xf767 */
            {8'h00}, /* 0xf766 */
            {8'h00}, /* 0xf765 */
            {8'h00}, /* 0xf764 */
            {8'h00}, /* 0xf763 */
            {8'h00}, /* 0xf762 */
            {8'h00}, /* 0xf761 */
            {8'h00}, /* 0xf760 */
            {8'h00}, /* 0xf75f */
            {8'h00}, /* 0xf75e */
            {8'h00}, /* 0xf75d */
            {8'h00}, /* 0xf75c */
            {8'h00}, /* 0xf75b */
            {8'h00}, /* 0xf75a */
            {8'h00}, /* 0xf759 */
            {8'h00}, /* 0xf758 */
            {8'h00}, /* 0xf757 */
            {8'h00}, /* 0xf756 */
            {8'h00}, /* 0xf755 */
            {8'h00}, /* 0xf754 */
            {8'h00}, /* 0xf753 */
            {8'h00}, /* 0xf752 */
            {8'h00}, /* 0xf751 */
            {8'h00}, /* 0xf750 */
            {8'h00}, /* 0xf74f */
            {8'h00}, /* 0xf74e */
            {8'h00}, /* 0xf74d */
            {8'h00}, /* 0xf74c */
            {8'h00}, /* 0xf74b */
            {8'h00}, /* 0xf74a */
            {8'h00}, /* 0xf749 */
            {8'h00}, /* 0xf748 */
            {8'h00}, /* 0xf747 */
            {8'h00}, /* 0xf746 */
            {8'h00}, /* 0xf745 */
            {8'h00}, /* 0xf744 */
            {8'h00}, /* 0xf743 */
            {8'h00}, /* 0xf742 */
            {8'h00}, /* 0xf741 */
            {8'h00}, /* 0xf740 */
            {8'h00}, /* 0xf73f */
            {8'h00}, /* 0xf73e */
            {8'h00}, /* 0xf73d */
            {8'h00}, /* 0xf73c */
            {8'h00}, /* 0xf73b */
            {8'h00}, /* 0xf73a */
            {8'h00}, /* 0xf739 */
            {8'h00}, /* 0xf738 */
            {8'h00}, /* 0xf737 */
            {8'h00}, /* 0xf736 */
            {8'h00}, /* 0xf735 */
            {8'h00}, /* 0xf734 */
            {8'h00}, /* 0xf733 */
            {8'h00}, /* 0xf732 */
            {8'h00}, /* 0xf731 */
            {8'h00}, /* 0xf730 */
            {8'h00}, /* 0xf72f */
            {8'h00}, /* 0xf72e */
            {8'h00}, /* 0xf72d */
            {8'h00}, /* 0xf72c */
            {8'h00}, /* 0xf72b */
            {8'h00}, /* 0xf72a */
            {8'h00}, /* 0xf729 */
            {8'h00}, /* 0xf728 */
            {8'h00}, /* 0xf727 */
            {8'h00}, /* 0xf726 */
            {8'h00}, /* 0xf725 */
            {8'h00}, /* 0xf724 */
            {8'h00}, /* 0xf723 */
            {8'h00}, /* 0xf722 */
            {8'h00}, /* 0xf721 */
            {8'h00}, /* 0xf720 */
            {8'h00}, /* 0xf71f */
            {8'h00}, /* 0xf71e */
            {8'h00}, /* 0xf71d */
            {8'h00}, /* 0xf71c */
            {8'h00}, /* 0xf71b */
            {8'h00}, /* 0xf71a */
            {8'h00}, /* 0xf719 */
            {8'h00}, /* 0xf718 */
            {8'h00}, /* 0xf717 */
            {8'h00}, /* 0xf716 */
            {8'h00}, /* 0xf715 */
            {8'h00}, /* 0xf714 */
            {8'h00}, /* 0xf713 */
            {8'h00}, /* 0xf712 */
            {8'h00}, /* 0xf711 */
            {8'h00}, /* 0xf710 */
            {8'h00}, /* 0xf70f */
            {8'h00}, /* 0xf70e */
            {8'h00}, /* 0xf70d */
            {8'h00}, /* 0xf70c */
            {8'h00}, /* 0xf70b */
            {8'h00}, /* 0xf70a */
            {8'h00}, /* 0xf709 */
            {8'h00}, /* 0xf708 */
            {8'h00}, /* 0xf707 */
            {8'h00}, /* 0xf706 */
            {8'h00}, /* 0xf705 */
            {8'h00}, /* 0xf704 */
            {8'h00}, /* 0xf703 */
            {8'h00}, /* 0xf702 */
            {8'h00}, /* 0xf701 */
            {8'h00}, /* 0xf700 */
            {8'h00}, /* 0xf6ff */
            {8'h00}, /* 0xf6fe */
            {8'h00}, /* 0xf6fd */
            {8'h00}, /* 0xf6fc */
            {8'h00}, /* 0xf6fb */
            {8'h00}, /* 0xf6fa */
            {8'h00}, /* 0xf6f9 */
            {8'h00}, /* 0xf6f8 */
            {8'h00}, /* 0xf6f7 */
            {8'h00}, /* 0xf6f6 */
            {8'h00}, /* 0xf6f5 */
            {8'h00}, /* 0xf6f4 */
            {8'h00}, /* 0xf6f3 */
            {8'h00}, /* 0xf6f2 */
            {8'h00}, /* 0xf6f1 */
            {8'h00}, /* 0xf6f0 */
            {8'h00}, /* 0xf6ef */
            {8'h00}, /* 0xf6ee */
            {8'h00}, /* 0xf6ed */
            {8'h00}, /* 0xf6ec */
            {8'h00}, /* 0xf6eb */
            {8'h00}, /* 0xf6ea */
            {8'h00}, /* 0xf6e9 */
            {8'h00}, /* 0xf6e8 */
            {8'h00}, /* 0xf6e7 */
            {8'h00}, /* 0xf6e6 */
            {8'h00}, /* 0xf6e5 */
            {8'h00}, /* 0xf6e4 */
            {8'h00}, /* 0xf6e3 */
            {8'h00}, /* 0xf6e2 */
            {8'h00}, /* 0xf6e1 */
            {8'h00}, /* 0xf6e0 */
            {8'h00}, /* 0xf6df */
            {8'h00}, /* 0xf6de */
            {8'h00}, /* 0xf6dd */
            {8'h00}, /* 0xf6dc */
            {8'h00}, /* 0xf6db */
            {8'h00}, /* 0xf6da */
            {8'h00}, /* 0xf6d9 */
            {8'h00}, /* 0xf6d8 */
            {8'h00}, /* 0xf6d7 */
            {8'h00}, /* 0xf6d6 */
            {8'h00}, /* 0xf6d5 */
            {8'h00}, /* 0xf6d4 */
            {8'h00}, /* 0xf6d3 */
            {8'h00}, /* 0xf6d2 */
            {8'h00}, /* 0xf6d1 */
            {8'h00}, /* 0xf6d0 */
            {8'h00}, /* 0xf6cf */
            {8'h00}, /* 0xf6ce */
            {8'h00}, /* 0xf6cd */
            {8'h00}, /* 0xf6cc */
            {8'h00}, /* 0xf6cb */
            {8'h00}, /* 0xf6ca */
            {8'h00}, /* 0xf6c9 */
            {8'h00}, /* 0xf6c8 */
            {8'h00}, /* 0xf6c7 */
            {8'h00}, /* 0xf6c6 */
            {8'h00}, /* 0xf6c5 */
            {8'h00}, /* 0xf6c4 */
            {8'h00}, /* 0xf6c3 */
            {8'h00}, /* 0xf6c2 */
            {8'h00}, /* 0xf6c1 */
            {8'h00}, /* 0xf6c0 */
            {8'h00}, /* 0xf6bf */
            {8'h00}, /* 0xf6be */
            {8'h00}, /* 0xf6bd */
            {8'h00}, /* 0xf6bc */
            {8'h00}, /* 0xf6bb */
            {8'h00}, /* 0xf6ba */
            {8'h00}, /* 0xf6b9 */
            {8'h00}, /* 0xf6b8 */
            {8'h00}, /* 0xf6b7 */
            {8'h00}, /* 0xf6b6 */
            {8'h00}, /* 0xf6b5 */
            {8'h00}, /* 0xf6b4 */
            {8'h00}, /* 0xf6b3 */
            {8'h00}, /* 0xf6b2 */
            {8'h00}, /* 0xf6b1 */
            {8'h00}, /* 0xf6b0 */
            {8'h00}, /* 0xf6af */
            {8'h00}, /* 0xf6ae */
            {8'h00}, /* 0xf6ad */
            {8'h00}, /* 0xf6ac */
            {8'h00}, /* 0xf6ab */
            {8'h00}, /* 0xf6aa */
            {8'h00}, /* 0xf6a9 */
            {8'h00}, /* 0xf6a8 */
            {8'h00}, /* 0xf6a7 */
            {8'h00}, /* 0xf6a6 */
            {8'h00}, /* 0xf6a5 */
            {8'h00}, /* 0xf6a4 */
            {8'h00}, /* 0xf6a3 */
            {8'h00}, /* 0xf6a2 */
            {8'h00}, /* 0xf6a1 */
            {8'h00}, /* 0xf6a0 */
            {8'h00}, /* 0xf69f */
            {8'h00}, /* 0xf69e */
            {8'h00}, /* 0xf69d */
            {8'h00}, /* 0xf69c */
            {8'h00}, /* 0xf69b */
            {8'h00}, /* 0xf69a */
            {8'h00}, /* 0xf699 */
            {8'h00}, /* 0xf698 */
            {8'h00}, /* 0xf697 */
            {8'h00}, /* 0xf696 */
            {8'h00}, /* 0xf695 */
            {8'h00}, /* 0xf694 */
            {8'h00}, /* 0xf693 */
            {8'h00}, /* 0xf692 */
            {8'h00}, /* 0xf691 */
            {8'h00}, /* 0xf690 */
            {8'h00}, /* 0xf68f */
            {8'h00}, /* 0xf68e */
            {8'h00}, /* 0xf68d */
            {8'h00}, /* 0xf68c */
            {8'h00}, /* 0xf68b */
            {8'h00}, /* 0xf68a */
            {8'h00}, /* 0xf689 */
            {8'h00}, /* 0xf688 */
            {8'h00}, /* 0xf687 */
            {8'h00}, /* 0xf686 */
            {8'h00}, /* 0xf685 */
            {8'h00}, /* 0xf684 */
            {8'h00}, /* 0xf683 */
            {8'h00}, /* 0xf682 */
            {8'h00}, /* 0xf681 */
            {8'h00}, /* 0xf680 */
            {8'h00}, /* 0xf67f */
            {8'h00}, /* 0xf67e */
            {8'h00}, /* 0xf67d */
            {8'h00}, /* 0xf67c */
            {8'h00}, /* 0xf67b */
            {8'h00}, /* 0xf67a */
            {8'h00}, /* 0xf679 */
            {8'h00}, /* 0xf678 */
            {8'h00}, /* 0xf677 */
            {8'h00}, /* 0xf676 */
            {8'h00}, /* 0xf675 */
            {8'h00}, /* 0xf674 */
            {8'h00}, /* 0xf673 */
            {8'h00}, /* 0xf672 */
            {8'h00}, /* 0xf671 */
            {8'h00}, /* 0xf670 */
            {8'h00}, /* 0xf66f */
            {8'h00}, /* 0xf66e */
            {8'h00}, /* 0xf66d */
            {8'h00}, /* 0xf66c */
            {8'h00}, /* 0xf66b */
            {8'h00}, /* 0xf66a */
            {8'h00}, /* 0xf669 */
            {8'h00}, /* 0xf668 */
            {8'h00}, /* 0xf667 */
            {8'h00}, /* 0xf666 */
            {8'h00}, /* 0xf665 */
            {8'h00}, /* 0xf664 */
            {8'h00}, /* 0xf663 */
            {8'h00}, /* 0xf662 */
            {8'h00}, /* 0xf661 */
            {8'h00}, /* 0xf660 */
            {8'h00}, /* 0xf65f */
            {8'h00}, /* 0xf65e */
            {8'h00}, /* 0xf65d */
            {8'h00}, /* 0xf65c */
            {8'h00}, /* 0xf65b */
            {8'h00}, /* 0xf65a */
            {8'h00}, /* 0xf659 */
            {8'h00}, /* 0xf658 */
            {8'h00}, /* 0xf657 */
            {8'h00}, /* 0xf656 */
            {8'h00}, /* 0xf655 */
            {8'h00}, /* 0xf654 */
            {8'h00}, /* 0xf653 */
            {8'h00}, /* 0xf652 */
            {8'h00}, /* 0xf651 */
            {8'h00}, /* 0xf650 */
            {8'h00}, /* 0xf64f */
            {8'h00}, /* 0xf64e */
            {8'h00}, /* 0xf64d */
            {8'h00}, /* 0xf64c */
            {8'h00}, /* 0xf64b */
            {8'h00}, /* 0xf64a */
            {8'h00}, /* 0xf649 */
            {8'h00}, /* 0xf648 */
            {8'h00}, /* 0xf647 */
            {8'h00}, /* 0xf646 */
            {8'h00}, /* 0xf645 */
            {8'h00}, /* 0xf644 */
            {8'h00}, /* 0xf643 */
            {8'h00}, /* 0xf642 */
            {8'h00}, /* 0xf641 */
            {8'h00}, /* 0xf640 */
            {8'h00}, /* 0xf63f */
            {8'h00}, /* 0xf63e */
            {8'h00}, /* 0xf63d */
            {8'h00}, /* 0xf63c */
            {8'h00}, /* 0xf63b */
            {8'h00}, /* 0xf63a */
            {8'h00}, /* 0xf639 */
            {8'h00}, /* 0xf638 */
            {8'h00}, /* 0xf637 */
            {8'h00}, /* 0xf636 */
            {8'h00}, /* 0xf635 */
            {8'h00}, /* 0xf634 */
            {8'h00}, /* 0xf633 */
            {8'h00}, /* 0xf632 */
            {8'h00}, /* 0xf631 */
            {8'h00}, /* 0xf630 */
            {8'h00}, /* 0xf62f */
            {8'h00}, /* 0xf62e */
            {8'h00}, /* 0xf62d */
            {8'h00}, /* 0xf62c */
            {8'h00}, /* 0xf62b */
            {8'h00}, /* 0xf62a */
            {8'h00}, /* 0xf629 */
            {8'h00}, /* 0xf628 */
            {8'h00}, /* 0xf627 */
            {8'h00}, /* 0xf626 */
            {8'h00}, /* 0xf625 */
            {8'h00}, /* 0xf624 */
            {8'h00}, /* 0xf623 */
            {8'h00}, /* 0xf622 */
            {8'h00}, /* 0xf621 */
            {8'h00}, /* 0xf620 */
            {8'h00}, /* 0xf61f */
            {8'h00}, /* 0xf61e */
            {8'h00}, /* 0xf61d */
            {8'h00}, /* 0xf61c */
            {8'h00}, /* 0xf61b */
            {8'h00}, /* 0xf61a */
            {8'h00}, /* 0xf619 */
            {8'h00}, /* 0xf618 */
            {8'h00}, /* 0xf617 */
            {8'h00}, /* 0xf616 */
            {8'h00}, /* 0xf615 */
            {8'h00}, /* 0xf614 */
            {8'h00}, /* 0xf613 */
            {8'h00}, /* 0xf612 */
            {8'h00}, /* 0xf611 */
            {8'h00}, /* 0xf610 */
            {8'h00}, /* 0xf60f */
            {8'h00}, /* 0xf60e */
            {8'h00}, /* 0xf60d */
            {8'h00}, /* 0xf60c */
            {8'h00}, /* 0xf60b */
            {8'h00}, /* 0xf60a */
            {8'h00}, /* 0xf609 */
            {8'h00}, /* 0xf608 */
            {8'h00}, /* 0xf607 */
            {8'h00}, /* 0xf606 */
            {8'h00}, /* 0xf605 */
            {8'h00}, /* 0xf604 */
            {8'h00}, /* 0xf603 */
            {8'h00}, /* 0xf602 */
            {8'h00}, /* 0xf601 */
            {8'h00}, /* 0xf600 */
            {8'h00}, /* 0xf5ff */
            {8'h00}, /* 0xf5fe */
            {8'h00}, /* 0xf5fd */
            {8'h00}, /* 0xf5fc */
            {8'h00}, /* 0xf5fb */
            {8'h00}, /* 0xf5fa */
            {8'h00}, /* 0xf5f9 */
            {8'h00}, /* 0xf5f8 */
            {8'h00}, /* 0xf5f7 */
            {8'h00}, /* 0xf5f6 */
            {8'h00}, /* 0xf5f5 */
            {8'h00}, /* 0xf5f4 */
            {8'h00}, /* 0xf5f3 */
            {8'h00}, /* 0xf5f2 */
            {8'h00}, /* 0xf5f1 */
            {8'h00}, /* 0xf5f0 */
            {8'h00}, /* 0xf5ef */
            {8'h00}, /* 0xf5ee */
            {8'h00}, /* 0xf5ed */
            {8'h00}, /* 0xf5ec */
            {8'h00}, /* 0xf5eb */
            {8'h00}, /* 0xf5ea */
            {8'h00}, /* 0xf5e9 */
            {8'h00}, /* 0xf5e8 */
            {8'h00}, /* 0xf5e7 */
            {8'h00}, /* 0xf5e6 */
            {8'h00}, /* 0xf5e5 */
            {8'h00}, /* 0xf5e4 */
            {8'h00}, /* 0xf5e3 */
            {8'h00}, /* 0xf5e2 */
            {8'h00}, /* 0xf5e1 */
            {8'h00}, /* 0xf5e0 */
            {8'h00}, /* 0xf5df */
            {8'h00}, /* 0xf5de */
            {8'h00}, /* 0xf5dd */
            {8'h00}, /* 0xf5dc */
            {8'h00}, /* 0xf5db */
            {8'h00}, /* 0xf5da */
            {8'h00}, /* 0xf5d9 */
            {8'h00}, /* 0xf5d8 */
            {8'h00}, /* 0xf5d7 */
            {8'h00}, /* 0xf5d6 */
            {8'h00}, /* 0xf5d5 */
            {8'h00}, /* 0xf5d4 */
            {8'h00}, /* 0xf5d3 */
            {8'h00}, /* 0xf5d2 */
            {8'h00}, /* 0xf5d1 */
            {8'h00}, /* 0xf5d0 */
            {8'h00}, /* 0xf5cf */
            {8'h00}, /* 0xf5ce */
            {8'h00}, /* 0xf5cd */
            {8'h00}, /* 0xf5cc */
            {8'h00}, /* 0xf5cb */
            {8'h00}, /* 0xf5ca */
            {8'h00}, /* 0xf5c9 */
            {8'h00}, /* 0xf5c8 */
            {8'h00}, /* 0xf5c7 */
            {8'h00}, /* 0xf5c6 */
            {8'h00}, /* 0xf5c5 */
            {8'h00}, /* 0xf5c4 */
            {8'h00}, /* 0xf5c3 */
            {8'h00}, /* 0xf5c2 */
            {8'h00}, /* 0xf5c1 */
            {8'h00}, /* 0xf5c0 */
            {8'h00}, /* 0xf5bf */
            {8'h00}, /* 0xf5be */
            {8'h00}, /* 0xf5bd */
            {8'h00}, /* 0xf5bc */
            {8'h00}, /* 0xf5bb */
            {8'h00}, /* 0xf5ba */
            {8'h00}, /* 0xf5b9 */
            {8'h00}, /* 0xf5b8 */
            {8'h00}, /* 0xf5b7 */
            {8'h00}, /* 0xf5b6 */
            {8'h00}, /* 0xf5b5 */
            {8'h00}, /* 0xf5b4 */
            {8'h00}, /* 0xf5b3 */
            {8'h00}, /* 0xf5b2 */
            {8'h00}, /* 0xf5b1 */
            {8'h00}, /* 0xf5b0 */
            {8'h00}, /* 0xf5af */
            {8'h00}, /* 0xf5ae */
            {8'h00}, /* 0xf5ad */
            {8'h00}, /* 0xf5ac */
            {8'h00}, /* 0xf5ab */
            {8'h00}, /* 0xf5aa */
            {8'h00}, /* 0xf5a9 */
            {8'h00}, /* 0xf5a8 */
            {8'h00}, /* 0xf5a7 */
            {8'h00}, /* 0xf5a6 */
            {8'h00}, /* 0xf5a5 */
            {8'h00}, /* 0xf5a4 */
            {8'h00}, /* 0xf5a3 */
            {8'h00}, /* 0xf5a2 */
            {8'h00}, /* 0xf5a1 */
            {8'h00}, /* 0xf5a0 */
            {8'h00}, /* 0xf59f */
            {8'h00}, /* 0xf59e */
            {8'h00}, /* 0xf59d */
            {8'h00}, /* 0xf59c */
            {8'h00}, /* 0xf59b */
            {8'h00}, /* 0xf59a */
            {8'h00}, /* 0xf599 */
            {8'h00}, /* 0xf598 */
            {8'h00}, /* 0xf597 */
            {8'h00}, /* 0xf596 */
            {8'h00}, /* 0xf595 */
            {8'h00}, /* 0xf594 */
            {8'h00}, /* 0xf593 */
            {8'h00}, /* 0xf592 */
            {8'h00}, /* 0xf591 */
            {8'h00}, /* 0xf590 */
            {8'h00}, /* 0xf58f */
            {8'h00}, /* 0xf58e */
            {8'h00}, /* 0xf58d */
            {8'h00}, /* 0xf58c */
            {8'h00}, /* 0xf58b */
            {8'h00}, /* 0xf58a */
            {8'h00}, /* 0xf589 */
            {8'h00}, /* 0xf588 */
            {8'h00}, /* 0xf587 */
            {8'h00}, /* 0xf586 */
            {8'h00}, /* 0xf585 */
            {8'h00}, /* 0xf584 */
            {8'h00}, /* 0xf583 */
            {8'h00}, /* 0xf582 */
            {8'h00}, /* 0xf581 */
            {8'h00}, /* 0xf580 */
            {8'h00}, /* 0xf57f */
            {8'h00}, /* 0xf57e */
            {8'h00}, /* 0xf57d */
            {8'h00}, /* 0xf57c */
            {8'h00}, /* 0xf57b */
            {8'h00}, /* 0xf57a */
            {8'h00}, /* 0xf579 */
            {8'h00}, /* 0xf578 */
            {8'h00}, /* 0xf577 */
            {8'h00}, /* 0xf576 */
            {8'h00}, /* 0xf575 */
            {8'h00}, /* 0xf574 */
            {8'h00}, /* 0xf573 */
            {8'h00}, /* 0xf572 */
            {8'h00}, /* 0xf571 */
            {8'h00}, /* 0xf570 */
            {8'h00}, /* 0xf56f */
            {8'h00}, /* 0xf56e */
            {8'h00}, /* 0xf56d */
            {8'h00}, /* 0xf56c */
            {8'h00}, /* 0xf56b */
            {8'h00}, /* 0xf56a */
            {8'h00}, /* 0xf569 */
            {8'h00}, /* 0xf568 */
            {8'h00}, /* 0xf567 */
            {8'h00}, /* 0xf566 */
            {8'h00}, /* 0xf565 */
            {8'h00}, /* 0xf564 */
            {8'h00}, /* 0xf563 */
            {8'h00}, /* 0xf562 */
            {8'h00}, /* 0xf561 */
            {8'h00}, /* 0xf560 */
            {8'h00}, /* 0xf55f */
            {8'h00}, /* 0xf55e */
            {8'h00}, /* 0xf55d */
            {8'h00}, /* 0xf55c */
            {8'h00}, /* 0xf55b */
            {8'h00}, /* 0xf55a */
            {8'h00}, /* 0xf559 */
            {8'h00}, /* 0xf558 */
            {8'h00}, /* 0xf557 */
            {8'h00}, /* 0xf556 */
            {8'h00}, /* 0xf555 */
            {8'h00}, /* 0xf554 */
            {8'h00}, /* 0xf553 */
            {8'h00}, /* 0xf552 */
            {8'h00}, /* 0xf551 */
            {8'h00}, /* 0xf550 */
            {8'h00}, /* 0xf54f */
            {8'h00}, /* 0xf54e */
            {8'h00}, /* 0xf54d */
            {8'h00}, /* 0xf54c */
            {8'h00}, /* 0xf54b */
            {8'h00}, /* 0xf54a */
            {8'h00}, /* 0xf549 */
            {8'h00}, /* 0xf548 */
            {8'h00}, /* 0xf547 */
            {8'h00}, /* 0xf546 */
            {8'h00}, /* 0xf545 */
            {8'h00}, /* 0xf544 */
            {8'h00}, /* 0xf543 */
            {8'h00}, /* 0xf542 */
            {8'h00}, /* 0xf541 */
            {8'h00}, /* 0xf540 */
            {8'h00}, /* 0xf53f */
            {8'h00}, /* 0xf53e */
            {8'h00}, /* 0xf53d */
            {8'h00}, /* 0xf53c */
            {8'h00}, /* 0xf53b */
            {8'h00}, /* 0xf53a */
            {8'h00}, /* 0xf539 */
            {8'h00}, /* 0xf538 */
            {8'h00}, /* 0xf537 */
            {8'h00}, /* 0xf536 */
            {8'h00}, /* 0xf535 */
            {8'h00}, /* 0xf534 */
            {8'h00}, /* 0xf533 */
            {8'h00}, /* 0xf532 */
            {8'h00}, /* 0xf531 */
            {8'h00}, /* 0xf530 */
            {8'h00}, /* 0xf52f */
            {8'h00}, /* 0xf52e */
            {8'h00}, /* 0xf52d */
            {8'h00}, /* 0xf52c */
            {8'h00}, /* 0xf52b */
            {8'h00}, /* 0xf52a */
            {8'h00}, /* 0xf529 */
            {8'h00}, /* 0xf528 */
            {8'h00}, /* 0xf527 */
            {8'h00}, /* 0xf526 */
            {8'h00}, /* 0xf525 */
            {8'h00}, /* 0xf524 */
            {8'h00}, /* 0xf523 */
            {8'h00}, /* 0xf522 */
            {8'h00}, /* 0xf521 */
            {8'h00}, /* 0xf520 */
            {8'h00}, /* 0xf51f */
            {8'h00}, /* 0xf51e */
            {8'h00}, /* 0xf51d */
            {8'h00}, /* 0xf51c */
            {8'h00}, /* 0xf51b */
            {8'h00}, /* 0xf51a */
            {8'h00}, /* 0xf519 */
            {8'h00}, /* 0xf518 */
            {8'h00}, /* 0xf517 */
            {8'h00}, /* 0xf516 */
            {8'h00}, /* 0xf515 */
            {8'h00}, /* 0xf514 */
            {8'h00}, /* 0xf513 */
            {8'h00}, /* 0xf512 */
            {8'h00}, /* 0xf511 */
            {8'h00}, /* 0xf510 */
            {8'h00}, /* 0xf50f */
            {8'h00}, /* 0xf50e */
            {8'h00}, /* 0xf50d */
            {8'h00}, /* 0xf50c */
            {8'h00}, /* 0xf50b */
            {8'h00}, /* 0xf50a */
            {8'h00}, /* 0xf509 */
            {8'h00}, /* 0xf508 */
            {8'h00}, /* 0xf507 */
            {8'h00}, /* 0xf506 */
            {8'h00}, /* 0xf505 */
            {8'h00}, /* 0xf504 */
            {8'h00}, /* 0xf503 */
            {8'h00}, /* 0xf502 */
            {8'h00}, /* 0xf501 */
            {8'h00}, /* 0xf500 */
            {8'h00}, /* 0xf4ff */
            {8'h00}, /* 0xf4fe */
            {8'h00}, /* 0xf4fd */
            {8'h00}, /* 0xf4fc */
            {8'h00}, /* 0xf4fb */
            {8'h00}, /* 0xf4fa */
            {8'h00}, /* 0xf4f9 */
            {8'h00}, /* 0xf4f8 */
            {8'h00}, /* 0xf4f7 */
            {8'h00}, /* 0xf4f6 */
            {8'h00}, /* 0xf4f5 */
            {8'h00}, /* 0xf4f4 */
            {8'h00}, /* 0xf4f3 */
            {8'h00}, /* 0xf4f2 */
            {8'h00}, /* 0xf4f1 */
            {8'h00}, /* 0xf4f0 */
            {8'h00}, /* 0xf4ef */
            {8'h00}, /* 0xf4ee */
            {8'h00}, /* 0xf4ed */
            {8'h00}, /* 0xf4ec */
            {8'h00}, /* 0xf4eb */
            {8'h00}, /* 0xf4ea */
            {8'h00}, /* 0xf4e9 */
            {8'h00}, /* 0xf4e8 */
            {8'h00}, /* 0xf4e7 */
            {8'h00}, /* 0xf4e6 */
            {8'h00}, /* 0xf4e5 */
            {8'h00}, /* 0xf4e4 */
            {8'h00}, /* 0xf4e3 */
            {8'h00}, /* 0xf4e2 */
            {8'h00}, /* 0xf4e1 */
            {8'h00}, /* 0xf4e0 */
            {8'h00}, /* 0xf4df */
            {8'h00}, /* 0xf4de */
            {8'h00}, /* 0xf4dd */
            {8'h00}, /* 0xf4dc */
            {8'h00}, /* 0xf4db */
            {8'h00}, /* 0xf4da */
            {8'h00}, /* 0xf4d9 */
            {8'h00}, /* 0xf4d8 */
            {8'h00}, /* 0xf4d7 */
            {8'h00}, /* 0xf4d6 */
            {8'h00}, /* 0xf4d5 */
            {8'h00}, /* 0xf4d4 */
            {8'h00}, /* 0xf4d3 */
            {8'h00}, /* 0xf4d2 */
            {8'h00}, /* 0xf4d1 */
            {8'h00}, /* 0xf4d0 */
            {8'h00}, /* 0xf4cf */
            {8'h00}, /* 0xf4ce */
            {8'h00}, /* 0xf4cd */
            {8'h00}, /* 0xf4cc */
            {8'h00}, /* 0xf4cb */
            {8'h00}, /* 0xf4ca */
            {8'h00}, /* 0xf4c9 */
            {8'h00}, /* 0xf4c8 */
            {8'h00}, /* 0xf4c7 */
            {8'h00}, /* 0xf4c6 */
            {8'h00}, /* 0xf4c5 */
            {8'h00}, /* 0xf4c4 */
            {8'h00}, /* 0xf4c3 */
            {8'h00}, /* 0xf4c2 */
            {8'h00}, /* 0xf4c1 */
            {8'h00}, /* 0xf4c0 */
            {8'h00}, /* 0xf4bf */
            {8'h00}, /* 0xf4be */
            {8'h00}, /* 0xf4bd */
            {8'h00}, /* 0xf4bc */
            {8'h00}, /* 0xf4bb */
            {8'h00}, /* 0xf4ba */
            {8'h00}, /* 0xf4b9 */
            {8'h00}, /* 0xf4b8 */
            {8'h00}, /* 0xf4b7 */
            {8'h00}, /* 0xf4b6 */
            {8'h00}, /* 0xf4b5 */
            {8'h00}, /* 0xf4b4 */
            {8'h00}, /* 0xf4b3 */
            {8'h00}, /* 0xf4b2 */
            {8'h00}, /* 0xf4b1 */
            {8'h00}, /* 0xf4b0 */
            {8'h00}, /* 0xf4af */
            {8'h00}, /* 0xf4ae */
            {8'h00}, /* 0xf4ad */
            {8'h00}, /* 0xf4ac */
            {8'h00}, /* 0xf4ab */
            {8'h00}, /* 0xf4aa */
            {8'h00}, /* 0xf4a9 */
            {8'h00}, /* 0xf4a8 */
            {8'h00}, /* 0xf4a7 */
            {8'h00}, /* 0xf4a6 */
            {8'h00}, /* 0xf4a5 */
            {8'h00}, /* 0xf4a4 */
            {8'h00}, /* 0xf4a3 */
            {8'h00}, /* 0xf4a2 */
            {8'h00}, /* 0xf4a1 */
            {8'h00}, /* 0xf4a0 */
            {8'h00}, /* 0xf49f */
            {8'h00}, /* 0xf49e */
            {8'h00}, /* 0xf49d */
            {8'h00}, /* 0xf49c */
            {8'h00}, /* 0xf49b */
            {8'h00}, /* 0xf49a */
            {8'h00}, /* 0xf499 */
            {8'h00}, /* 0xf498 */
            {8'h00}, /* 0xf497 */
            {8'h00}, /* 0xf496 */
            {8'h00}, /* 0xf495 */
            {8'h00}, /* 0xf494 */
            {8'h00}, /* 0xf493 */
            {8'h00}, /* 0xf492 */
            {8'h00}, /* 0xf491 */
            {8'h00}, /* 0xf490 */
            {8'h00}, /* 0xf48f */
            {8'h00}, /* 0xf48e */
            {8'h00}, /* 0xf48d */
            {8'h00}, /* 0xf48c */
            {8'h00}, /* 0xf48b */
            {8'h00}, /* 0xf48a */
            {8'h00}, /* 0xf489 */
            {8'h00}, /* 0xf488 */
            {8'h00}, /* 0xf487 */
            {8'h00}, /* 0xf486 */
            {8'h00}, /* 0xf485 */
            {8'h00}, /* 0xf484 */
            {8'h00}, /* 0xf483 */
            {8'h00}, /* 0xf482 */
            {8'h00}, /* 0xf481 */
            {8'h00}, /* 0xf480 */
            {8'h00}, /* 0xf47f */
            {8'h00}, /* 0xf47e */
            {8'h00}, /* 0xf47d */
            {8'h00}, /* 0xf47c */
            {8'h00}, /* 0xf47b */
            {8'h00}, /* 0xf47a */
            {8'h00}, /* 0xf479 */
            {8'h00}, /* 0xf478 */
            {8'h00}, /* 0xf477 */
            {8'h00}, /* 0xf476 */
            {8'h00}, /* 0xf475 */
            {8'h00}, /* 0xf474 */
            {8'h00}, /* 0xf473 */
            {8'h00}, /* 0xf472 */
            {8'h00}, /* 0xf471 */
            {8'h00}, /* 0xf470 */
            {8'h00}, /* 0xf46f */
            {8'h00}, /* 0xf46e */
            {8'h00}, /* 0xf46d */
            {8'h00}, /* 0xf46c */
            {8'h00}, /* 0xf46b */
            {8'h00}, /* 0xf46a */
            {8'h00}, /* 0xf469 */
            {8'h00}, /* 0xf468 */
            {8'h00}, /* 0xf467 */
            {8'h00}, /* 0xf466 */
            {8'h00}, /* 0xf465 */
            {8'h00}, /* 0xf464 */
            {8'h00}, /* 0xf463 */
            {8'h00}, /* 0xf462 */
            {8'h00}, /* 0xf461 */
            {8'h00}, /* 0xf460 */
            {8'h00}, /* 0xf45f */
            {8'h00}, /* 0xf45e */
            {8'h00}, /* 0xf45d */
            {8'h00}, /* 0xf45c */
            {8'h00}, /* 0xf45b */
            {8'h00}, /* 0xf45a */
            {8'h00}, /* 0xf459 */
            {8'h00}, /* 0xf458 */
            {8'h00}, /* 0xf457 */
            {8'h00}, /* 0xf456 */
            {8'h00}, /* 0xf455 */
            {8'h00}, /* 0xf454 */
            {8'h00}, /* 0xf453 */
            {8'h00}, /* 0xf452 */
            {8'h00}, /* 0xf451 */
            {8'h00}, /* 0xf450 */
            {8'h00}, /* 0xf44f */
            {8'h00}, /* 0xf44e */
            {8'h00}, /* 0xf44d */
            {8'h00}, /* 0xf44c */
            {8'h00}, /* 0xf44b */
            {8'h00}, /* 0xf44a */
            {8'h00}, /* 0xf449 */
            {8'h00}, /* 0xf448 */
            {8'h00}, /* 0xf447 */
            {8'h00}, /* 0xf446 */
            {8'h00}, /* 0xf445 */
            {8'h00}, /* 0xf444 */
            {8'h00}, /* 0xf443 */
            {8'h00}, /* 0xf442 */
            {8'h00}, /* 0xf441 */
            {8'h00}, /* 0xf440 */
            {8'h00}, /* 0xf43f */
            {8'h00}, /* 0xf43e */
            {8'h00}, /* 0xf43d */
            {8'h00}, /* 0xf43c */
            {8'h00}, /* 0xf43b */
            {8'h00}, /* 0xf43a */
            {8'h00}, /* 0xf439 */
            {8'h00}, /* 0xf438 */
            {8'h00}, /* 0xf437 */
            {8'h00}, /* 0xf436 */
            {8'h00}, /* 0xf435 */
            {8'h00}, /* 0xf434 */
            {8'h00}, /* 0xf433 */
            {8'h00}, /* 0xf432 */
            {8'h00}, /* 0xf431 */
            {8'h00}, /* 0xf430 */
            {8'h00}, /* 0xf42f */
            {8'h00}, /* 0xf42e */
            {8'h00}, /* 0xf42d */
            {8'h00}, /* 0xf42c */
            {8'h00}, /* 0xf42b */
            {8'h00}, /* 0xf42a */
            {8'h00}, /* 0xf429 */
            {8'h00}, /* 0xf428 */
            {8'h00}, /* 0xf427 */
            {8'h00}, /* 0xf426 */
            {8'h00}, /* 0xf425 */
            {8'h00}, /* 0xf424 */
            {8'h00}, /* 0xf423 */
            {8'h00}, /* 0xf422 */
            {8'h00}, /* 0xf421 */
            {8'h00}, /* 0xf420 */
            {8'h00}, /* 0xf41f */
            {8'h00}, /* 0xf41e */
            {8'h00}, /* 0xf41d */
            {8'h00}, /* 0xf41c */
            {8'h00}, /* 0xf41b */
            {8'h00}, /* 0xf41a */
            {8'h00}, /* 0xf419 */
            {8'h00}, /* 0xf418 */
            {8'h00}, /* 0xf417 */
            {8'h00}, /* 0xf416 */
            {8'h00}, /* 0xf415 */
            {8'h00}, /* 0xf414 */
            {8'h00}, /* 0xf413 */
            {8'h00}, /* 0xf412 */
            {8'h00}, /* 0xf411 */
            {8'h00}, /* 0xf410 */
            {8'h00}, /* 0xf40f */
            {8'h00}, /* 0xf40e */
            {8'h00}, /* 0xf40d */
            {8'h00}, /* 0xf40c */
            {8'h00}, /* 0xf40b */
            {8'h00}, /* 0xf40a */
            {8'h00}, /* 0xf409 */
            {8'h00}, /* 0xf408 */
            {8'h00}, /* 0xf407 */
            {8'h00}, /* 0xf406 */
            {8'h00}, /* 0xf405 */
            {8'h00}, /* 0xf404 */
            {8'h00}, /* 0xf403 */
            {8'h00}, /* 0xf402 */
            {8'h00}, /* 0xf401 */
            {8'h00}, /* 0xf400 */
            {8'h00}, /* 0xf3ff */
            {8'h00}, /* 0xf3fe */
            {8'h00}, /* 0xf3fd */
            {8'h00}, /* 0xf3fc */
            {8'h00}, /* 0xf3fb */
            {8'h00}, /* 0xf3fa */
            {8'h00}, /* 0xf3f9 */
            {8'h00}, /* 0xf3f8 */
            {8'h00}, /* 0xf3f7 */
            {8'h00}, /* 0xf3f6 */
            {8'h00}, /* 0xf3f5 */
            {8'h00}, /* 0xf3f4 */
            {8'h00}, /* 0xf3f3 */
            {8'h00}, /* 0xf3f2 */
            {8'h00}, /* 0xf3f1 */
            {8'h00}, /* 0xf3f0 */
            {8'h00}, /* 0xf3ef */
            {8'h00}, /* 0xf3ee */
            {8'h00}, /* 0xf3ed */
            {8'h00}, /* 0xf3ec */
            {8'h00}, /* 0xf3eb */
            {8'h00}, /* 0xf3ea */
            {8'h00}, /* 0xf3e9 */
            {8'h00}, /* 0xf3e8 */
            {8'h00}, /* 0xf3e7 */
            {8'h00}, /* 0xf3e6 */
            {8'h00}, /* 0xf3e5 */
            {8'h00}, /* 0xf3e4 */
            {8'h00}, /* 0xf3e3 */
            {8'h00}, /* 0xf3e2 */
            {8'h00}, /* 0xf3e1 */
            {8'h00}, /* 0xf3e0 */
            {8'h00}, /* 0xf3df */
            {8'h00}, /* 0xf3de */
            {8'h00}, /* 0xf3dd */
            {8'h00}, /* 0xf3dc */
            {8'h00}, /* 0xf3db */
            {8'h00}, /* 0xf3da */
            {8'h00}, /* 0xf3d9 */
            {8'h00}, /* 0xf3d8 */
            {8'h00}, /* 0xf3d7 */
            {8'h00}, /* 0xf3d6 */
            {8'h00}, /* 0xf3d5 */
            {8'h00}, /* 0xf3d4 */
            {8'h00}, /* 0xf3d3 */
            {8'h00}, /* 0xf3d2 */
            {8'h00}, /* 0xf3d1 */
            {8'h00}, /* 0xf3d0 */
            {8'h00}, /* 0xf3cf */
            {8'h00}, /* 0xf3ce */
            {8'h00}, /* 0xf3cd */
            {8'h00}, /* 0xf3cc */
            {8'h00}, /* 0xf3cb */
            {8'h00}, /* 0xf3ca */
            {8'h00}, /* 0xf3c9 */
            {8'h00}, /* 0xf3c8 */
            {8'h00}, /* 0xf3c7 */
            {8'h00}, /* 0xf3c6 */
            {8'h00}, /* 0xf3c5 */
            {8'h00}, /* 0xf3c4 */
            {8'h00}, /* 0xf3c3 */
            {8'h00}, /* 0xf3c2 */
            {8'h00}, /* 0xf3c1 */
            {8'h00}, /* 0xf3c0 */
            {8'h00}, /* 0xf3bf */
            {8'h00}, /* 0xf3be */
            {8'h00}, /* 0xf3bd */
            {8'h00}, /* 0xf3bc */
            {8'h00}, /* 0xf3bb */
            {8'h00}, /* 0xf3ba */
            {8'h00}, /* 0xf3b9 */
            {8'h00}, /* 0xf3b8 */
            {8'h00}, /* 0xf3b7 */
            {8'h00}, /* 0xf3b6 */
            {8'h00}, /* 0xf3b5 */
            {8'h00}, /* 0xf3b4 */
            {8'h00}, /* 0xf3b3 */
            {8'h00}, /* 0xf3b2 */
            {8'h00}, /* 0xf3b1 */
            {8'h00}, /* 0xf3b0 */
            {8'h00}, /* 0xf3af */
            {8'h00}, /* 0xf3ae */
            {8'h00}, /* 0xf3ad */
            {8'h00}, /* 0xf3ac */
            {8'h00}, /* 0xf3ab */
            {8'h00}, /* 0xf3aa */
            {8'h00}, /* 0xf3a9 */
            {8'h00}, /* 0xf3a8 */
            {8'h00}, /* 0xf3a7 */
            {8'h00}, /* 0xf3a6 */
            {8'h00}, /* 0xf3a5 */
            {8'h00}, /* 0xf3a4 */
            {8'h00}, /* 0xf3a3 */
            {8'h00}, /* 0xf3a2 */
            {8'h00}, /* 0xf3a1 */
            {8'h00}, /* 0xf3a0 */
            {8'h00}, /* 0xf39f */
            {8'h00}, /* 0xf39e */
            {8'h00}, /* 0xf39d */
            {8'h00}, /* 0xf39c */
            {8'h00}, /* 0xf39b */
            {8'h00}, /* 0xf39a */
            {8'h00}, /* 0xf399 */
            {8'h00}, /* 0xf398 */
            {8'h00}, /* 0xf397 */
            {8'h00}, /* 0xf396 */
            {8'h00}, /* 0xf395 */
            {8'h00}, /* 0xf394 */
            {8'h00}, /* 0xf393 */
            {8'h00}, /* 0xf392 */
            {8'h00}, /* 0xf391 */
            {8'h00}, /* 0xf390 */
            {8'h00}, /* 0xf38f */
            {8'h00}, /* 0xf38e */
            {8'h00}, /* 0xf38d */
            {8'h00}, /* 0xf38c */
            {8'h00}, /* 0xf38b */
            {8'h00}, /* 0xf38a */
            {8'h00}, /* 0xf389 */
            {8'h00}, /* 0xf388 */
            {8'h00}, /* 0xf387 */
            {8'h00}, /* 0xf386 */
            {8'h00}, /* 0xf385 */
            {8'h00}, /* 0xf384 */
            {8'h00}, /* 0xf383 */
            {8'h00}, /* 0xf382 */
            {8'h00}, /* 0xf381 */
            {8'h00}, /* 0xf380 */
            {8'h00}, /* 0xf37f */
            {8'h00}, /* 0xf37e */
            {8'h00}, /* 0xf37d */
            {8'h00}, /* 0xf37c */
            {8'h00}, /* 0xf37b */
            {8'h00}, /* 0xf37a */
            {8'h00}, /* 0xf379 */
            {8'h00}, /* 0xf378 */
            {8'h00}, /* 0xf377 */
            {8'h00}, /* 0xf376 */
            {8'h00}, /* 0xf375 */
            {8'h00}, /* 0xf374 */
            {8'h00}, /* 0xf373 */
            {8'h00}, /* 0xf372 */
            {8'h00}, /* 0xf371 */
            {8'h00}, /* 0xf370 */
            {8'h00}, /* 0xf36f */
            {8'h00}, /* 0xf36e */
            {8'h00}, /* 0xf36d */
            {8'h00}, /* 0xf36c */
            {8'h00}, /* 0xf36b */
            {8'h00}, /* 0xf36a */
            {8'h00}, /* 0xf369 */
            {8'h00}, /* 0xf368 */
            {8'h00}, /* 0xf367 */
            {8'h00}, /* 0xf366 */
            {8'h00}, /* 0xf365 */
            {8'h00}, /* 0xf364 */
            {8'h00}, /* 0xf363 */
            {8'h00}, /* 0xf362 */
            {8'h00}, /* 0xf361 */
            {8'h00}, /* 0xf360 */
            {8'h00}, /* 0xf35f */
            {8'h00}, /* 0xf35e */
            {8'h00}, /* 0xf35d */
            {8'h00}, /* 0xf35c */
            {8'h00}, /* 0xf35b */
            {8'h00}, /* 0xf35a */
            {8'h00}, /* 0xf359 */
            {8'h00}, /* 0xf358 */
            {8'h00}, /* 0xf357 */
            {8'h00}, /* 0xf356 */
            {8'h00}, /* 0xf355 */
            {8'h00}, /* 0xf354 */
            {8'h00}, /* 0xf353 */
            {8'h00}, /* 0xf352 */
            {8'h00}, /* 0xf351 */
            {8'h00}, /* 0xf350 */
            {8'h00}, /* 0xf34f */
            {8'h00}, /* 0xf34e */
            {8'h00}, /* 0xf34d */
            {8'h00}, /* 0xf34c */
            {8'h00}, /* 0xf34b */
            {8'h00}, /* 0xf34a */
            {8'h00}, /* 0xf349 */
            {8'h00}, /* 0xf348 */
            {8'h00}, /* 0xf347 */
            {8'h00}, /* 0xf346 */
            {8'h00}, /* 0xf345 */
            {8'h00}, /* 0xf344 */
            {8'h00}, /* 0xf343 */
            {8'h00}, /* 0xf342 */
            {8'h00}, /* 0xf341 */
            {8'h00}, /* 0xf340 */
            {8'h00}, /* 0xf33f */
            {8'h00}, /* 0xf33e */
            {8'h00}, /* 0xf33d */
            {8'h00}, /* 0xf33c */
            {8'h00}, /* 0xf33b */
            {8'h00}, /* 0xf33a */
            {8'h00}, /* 0xf339 */
            {8'h00}, /* 0xf338 */
            {8'h00}, /* 0xf337 */
            {8'h00}, /* 0xf336 */
            {8'h00}, /* 0xf335 */
            {8'h00}, /* 0xf334 */
            {8'h00}, /* 0xf333 */
            {8'h00}, /* 0xf332 */
            {8'h00}, /* 0xf331 */
            {8'h00}, /* 0xf330 */
            {8'h00}, /* 0xf32f */
            {8'h00}, /* 0xf32e */
            {8'h00}, /* 0xf32d */
            {8'h00}, /* 0xf32c */
            {8'h00}, /* 0xf32b */
            {8'h00}, /* 0xf32a */
            {8'h00}, /* 0xf329 */
            {8'h00}, /* 0xf328 */
            {8'h00}, /* 0xf327 */
            {8'h00}, /* 0xf326 */
            {8'h00}, /* 0xf325 */
            {8'h00}, /* 0xf324 */
            {8'h00}, /* 0xf323 */
            {8'h00}, /* 0xf322 */
            {8'h00}, /* 0xf321 */
            {8'h00}, /* 0xf320 */
            {8'h00}, /* 0xf31f */
            {8'h00}, /* 0xf31e */
            {8'h00}, /* 0xf31d */
            {8'h00}, /* 0xf31c */
            {8'h00}, /* 0xf31b */
            {8'h00}, /* 0xf31a */
            {8'h00}, /* 0xf319 */
            {8'h00}, /* 0xf318 */
            {8'h00}, /* 0xf317 */
            {8'h00}, /* 0xf316 */
            {8'h00}, /* 0xf315 */
            {8'h00}, /* 0xf314 */
            {8'h00}, /* 0xf313 */
            {8'h00}, /* 0xf312 */
            {8'h00}, /* 0xf311 */
            {8'h00}, /* 0xf310 */
            {8'h00}, /* 0xf30f */
            {8'h00}, /* 0xf30e */
            {8'h00}, /* 0xf30d */
            {8'h00}, /* 0xf30c */
            {8'h00}, /* 0xf30b */
            {8'h00}, /* 0xf30a */
            {8'h00}, /* 0xf309 */
            {8'h00}, /* 0xf308 */
            {8'h00}, /* 0xf307 */
            {8'h00}, /* 0xf306 */
            {8'h00}, /* 0xf305 */
            {8'h00}, /* 0xf304 */
            {8'h00}, /* 0xf303 */
            {8'h00}, /* 0xf302 */
            {8'h00}, /* 0xf301 */
            {8'h00}, /* 0xf300 */
            {8'h00}, /* 0xf2ff */
            {8'h00}, /* 0xf2fe */
            {8'h00}, /* 0xf2fd */
            {8'h00}, /* 0xf2fc */
            {8'h00}, /* 0xf2fb */
            {8'h00}, /* 0xf2fa */
            {8'h00}, /* 0xf2f9 */
            {8'h00}, /* 0xf2f8 */
            {8'h00}, /* 0xf2f7 */
            {8'h00}, /* 0xf2f6 */
            {8'h00}, /* 0xf2f5 */
            {8'h00}, /* 0xf2f4 */
            {8'h00}, /* 0xf2f3 */
            {8'h00}, /* 0xf2f2 */
            {8'h00}, /* 0xf2f1 */
            {8'h00}, /* 0xf2f0 */
            {8'h00}, /* 0xf2ef */
            {8'h00}, /* 0xf2ee */
            {8'h00}, /* 0xf2ed */
            {8'h00}, /* 0xf2ec */
            {8'h00}, /* 0xf2eb */
            {8'h00}, /* 0xf2ea */
            {8'h00}, /* 0xf2e9 */
            {8'h00}, /* 0xf2e8 */
            {8'h00}, /* 0xf2e7 */
            {8'h00}, /* 0xf2e6 */
            {8'h00}, /* 0xf2e5 */
            {8'h00}, /* 0xf2e4 */
            {8'h00}, /* 0xf2e3 */
            {8'h00}, /* 0xf2e2 */
            {8'h00}, /* 0xf2e1 */
            {8'h00}, /* 0xf2e0 */
            {8'h00}, /* 0xf2df */
            {8'h00}, /* 0xf2de */
            {8'h00}, /* 0xf2dd */
            {8'h00}, /* 0xf2dc */
            {8'h00}, /* 0xf2db */
            {8'h00}, /* 0xf2da */
            {8'h00}, /* 0xf2d9 */
            {8'h00}, /* 0xf2d8 */
            {8'h00}, /* 0xf2d7 */
            {8'h00}, /* 0xf2d6 */
            {8'h00}, /* 0xf2d5 */
            {8'h00}, /* 0xf2d4 */
            {8'h00}, /* 0xf2d3 */
            {8'h00}, /* 0xf2d2 */
            {8'h00}, /* 0xf2d1 */
            {8'h00}, /* 0xf2d0 */
            {8'h00}, /* 0xf2cf */
            {8'h00}, /* 0xf2ce */
            {8'h00}, /* 0xf2cd */
            {8'h00}, /* 0xf2cc */
            {8'h00}, /* 0xf2cb */
            {8'h00}, /* 0xf2ca */
            {8'h00}, /* 0xf2c9 */
            {8'h00}, /* 0xf2c8 */
            {8'h00}, /* 0xf2c7 */
            {8'h00}, /* 0xf2c6 */
            {8'h00}, /* 0xf2c5 */
            {8'h00}, /* 0xf2c4 */
            {8'h00}, /* 0xf2c3 */
            {8'h00}, /* 0xf2c2 */
            {8'h00}, /* 0xf2c1 */
            {8'h00}, /* 0xf2c0 */
            {8'h00}, /* 0xf2bf */
            {8'h00}, /* 0xf2be */
            {8'h00}, /* 0xf2bd */
            {8'h00}, /* 0xf2bc */
            {8'h00}, /* 0xf2bb */
            {8'h00}, /* 0xf2ba */
            {8'h00}, /* 0xf2b9 */
            {8'h00}, /* 0xf2b8 */
            {8'h00}, /* 0xf2b7 */
            {8'h00}, /* 0xf2b6 */
            {8'h00}, /* 0xf2b5 */
            {8'h00}, /* 0xf2b4 */
            {8'h00}, /* 0xf2b3 */
            {8'h00}, /* 0xf2b2 */
            {8'h00}, /* 0xf2b1 */
            {8'h00}, /* 0xf2b0 */
            {8'h00}, /* 0xf2af */
            {8'h00}, /* 0xf2ae */
            {8'h00}, /* 0xf2ad */
            {8'h00}, /* 0xf2ac */
            {8'h00}, /* 0xf2ab */
            {8'h00}, /* 0xf2aa */
            {8'h00}, /* 0xf2a9 */
            {8'h00}, /* 0xf2a8 */
            {8'h00}, /* 0xf2a7 */
            {8'h00}, /* 0xf2a6 */
            {8'h00}, /* 0xf2a5 */
            {8'h00}, /* 0xf2a4 */
            {8'h00}, /* 0xf2a3 */
            {8'h00}, /* 0xf2a2 */
            {8'h00}, /* 0xf2a1 */
            {8'h00}, /* 0xf2a0 */
            {8'h00}, /* 0xf29f */
            {8'h00}, /* 0xf29e */
            {8'h00}, /* 0xf29d */
            {8'h00}, /* 0xf29c */
            {8'h00}, /* 0xf29b */
            {8'h00}, /* 0xf29a */
            {8'h00}, /* 0xf299 */
            {8'h00}, /* 0xf298 */
            {8'h00}, /* 0xf297 */
            {8'h00}, /* 0xf296 */
            {8'h00}, /* 0xf295 */
            {8'h00}, /* 0xf294 */
            {8'h00}, /* 0xf293 */
            {8'h00}, /* 0xf292 */
            {8'h00}, /* 0xf291 */
            {8'h00}, /* 0xf290 */
            {8'h00}, /* 0xf28f */
            {8'h00}, /* 0xf28e */
            {8'h00}, /* 0xf28d */
            {8'h00}, /* 0xf28c */
            {8'h00}, /* 0xf28b */
            {8'h00}, /* 0xf28a */
            {8'h00}, /* 0xf289 */
            {8'h00}, /* 0xf288 */
            {8'h00}, /* 0xf287 */
            {8'h00}, /* 0xf286 */
            {8'h00}, /* 0xf285 */
            {8'h00}, /* 0xf284 */
            {8'h00}, /* 0xf283 */
            {8'h00}, /* 0xf282 */
            {8'h00}, /* 0xf281 */
            {8'h00}, /* 0xf280 */
            {8'h00}, /* 0xf27f */
            {8'h00}, /* 0xf27e */
            {8'h00}, /* 0xf27d */
            {8'h00}, /* 0xf27c */
            {8'h00}, /* 0xf27b */
            {8'h00}, /* 0xf27a */
            {8'h00}, /* 0xf279 */
            {8'h00}, /* 0xf278 */
            {8'h00}, /* 0xf277 */
            {8'h00}, /* 0xf276 */
            {8'h00}, /* 0xf275 */
            {8'h00}, /* 0xf274 */
            {8'h00}, /* 0xf273 */
            {8'h00}, /* 0xf272 */
            {8'h00}, /* 0xf271 */
            {8'h00}, /* 0xf270 */
            {8'h00}, /* 0xf26f */
            {8'h00}, /* 0xf26e */
            {8'h00}, /* 0xf26d */
            {8'h00}, /* 0xf26c */
            {8'h00}, /* 0xf26b */
            {8'h00}, /* 0xf26a */
            {8'h00}, /* 0xf269 */
            {8'h00}, /* 0xf268 */
            {8'h00}, /* 0xf267 */
            {8'h00}, /* 0xf266 */
            {8'h00}, /* 0xf265 */
            {8'h00}, /* 0xf264 */
            {8'h00}, /* 0xf263 */
            {8'h00}, /* 0xf262 */
            {8'h00}, /* 0xf261 */
            {8'h00}, /* 0xf260 */
            {8'h00}, /* 0xf25f */
            {8'h00}, /* 0xf25e */
            {8'h00}, /* 0xf25d */
            {8'h00}, /* 0xf25c */
            {8'h00}, /* 0xf25b */
            {8'h00}, /* 0xf25a */
            {8'h00}, /* 0xf259 */
            {8'h00}, /* 0xf258 */
            {8'h00}, /* 0xf257 */
            {8'h00}, /* 0xf256 */
            {8'h00}, /* 0xf255 */
            {8'h00}, /* 0xf254 */
            {8'h00}, /* 0xf253 */
            {8'h00}, /* 0xf252 */
            {8'h00}, /* 0xf251 */
            {8'h00}, /* 0xf250 */
            {8'h00}, /* 0xf24f */
            {8'h00}, /* 0xf24e */
            {8'h00}, /* 0xf24d */
            {8'h00}, /* 0xf24c */
            {8'h00}, /* 0xf24b */
            {8'h00}, /* 0xf24a */
            {8'h00}, /* 0xf249 */
            {8'h00}, /* 0xf248 */
            {8'h00}, /* 0xf247 */
            {8'h00}, /* 0xf246 */
            {8'h00}, /* 0xf245 */
            {8'h00}, /* 0xf244 */
            {8'h00}, /* 0xf243 */
            {8'h00}, /* 0xf242 */
            {8'h00}, /* 0xf241 */
            {8'h00}, /* 0xf240 */
            {8'h00}, /* 0xf23f */
            {8'h00}, /* 0xf23e */
            {8'h00}, /* 0xf23d */
            {8'h00}, /* 0xf23c */
            {8'h00}, /* 0xf23b */
            {8'h00}, /* 0xf23a */
            {8'h00}, /* 0xf239 */
            {8'h00}, /* 0xf238 */
            {8'h00}, /* 0xf237 */
            {8'h00}, /* 0xf236 */
            {8'h00}, /* 0xf235 */
            {8'h00}, /* 0xf234 */
            {8'h00}, /* 0xf233 */
            {8'h00}, /* 0xf232 */
            {8'h00}, /* 0xf231 */
            {8'h00}, /* 0xf230 */
            {8'h00}, /* 0xf22f */
            {8'h00}, /* 0xf22e */
            {8'h00}, /* 0xf22d */
            {8'h00}, /* 0xf22c */
            {8'h00}, /* 0xf22b */
            {8'h00}, /* 0xf22a */
            {8'h00}, /* 0xf229 */
            {8'h00}, /* 0xf228 */
            {8'h00}, /* 0xf227 */
            {8'h00}, /* 0xf226 */
            {8'h00}, /* 0xf225 */
            {8'h00}, /* 0xf224 */
            {8'h00}, /* 0xf223 */
            {8'h00}, /* 0xf222 */
            {8'h00}, /* 0xf221 */
            {8'h00}, /* 0xf220 */
            {8'h00}, /* 0xf21f */
            {8'h00}, /* 0xf21e */
            {8'h00}, /* 0xf21d */
            {8'h00}, /* 0xf21c */
            {8'h00}, /* 0xf21b */
            {8'h00}, /* 0xf21a */
            {8'h00}, /* 0xf219 */
            {8'h00}, /* 0xf218 */
            {8'h00}, /* 0xf217 */
            {8'h00}, /* 0xf216 */
            {8'h00}, /* 0xf215 */
            {8'h00}, /* 0xf214 */
            {8'h00}, /* 0xf213 */
            {8'h00}, /* 0xf212 */
            {8'h00}, /* 0xf211 */
            {8'h00}, /* 0xf210 */
            {8'h00}, /* 0xf20f */
            {8'h00}, /* 0xf20e */
            {8'h00}, /* 0xf20d */
            {8'h00}, /* 0xf20c */
            {8'h00}, /* 0xf20b */
            {8'h00}, /* 0xf20a */
            {8'h00}, /* 0xf209 */
            {8'h00}, /* 0xf208 */
            {8'h00}, /* 0xf207 */
            {8'h00}, /* 0xf206 */
            {8'h00}, /* 0xf205 */
            {8'h00}, /* 0xf204 */
            {8'h00}, /* 0xf203 */
            {8'h00}, /* 0xf202 */
            {8'h00}, /* 0xf201 */
            {8'h00}, /* 0xf200 */
            {8'h00}, /* 0xf1ff */
            {8'h00}, /* 0xf1fe */
            {8'h00}, /* 0xf1fd */
            {8'h00}, /* 0xf1fc */
            {8'h00}, /* 0xf1fb */
            {8'h00}, /* 0xf1fa */
            {8'h00}, /* 0xf1f9 */
            {8'h00}, /* 0xf1f8 */
            {8'h00}, /* 0xf1f7 */
            {8'h00}, /* 0xf1f6 */
            {8'h00}, /* 0xf1f5 */
            {8'h00}, /* 0xf1f4 */
            {8'h00}, /* 0xf1f3 */
            {8'h00}, /* 0xf1f2 */
            {8'h00}, /* 0xf1f1 */
            {8'h00}, /* 0xf1f0 */
            {8'h00}, /* 0xf1ef */
            {8'h00}, /* 0xf1ee */
            {8'h00}, /* 0xf1ed */
            {8'h00}, /* 0xf1ec */
            {8'h00}, /* 0xf1eb */
            {8'h00}, /* 0xf1ea */
            {8'h00}, /* 0xf1e9 */
            {8'h00}, /* 0xf1e8 */
            {8'h00}, /* 0xf1e7 */
            {8'h00}, /* 0xf1e6 */
            {8'h00}, /* 0xf1e5 */
            {8'h00}, /* 0xf1e4 */
            {8'h00}, /* 0xf1e3 */
            {8'h00}, /* 0xf1e2 */
            {8'h00}, /* 0xf1e1 */
            {8'h00}, /* 0xf1e0 */
            {8'h00}, /* 0xf1df */
            {8'h00}, /* 0xf1de */
            {8'h00}, /* 0xf1dd */
            {8'h00}, /* 0xf1dc */
            {8'h00}, /* 0xf1db */
            {8'h00}, /* 0xf1da */
            {8'h00}, /* 0xf1d9 */
            {8'h00}, /* 0xf1d8 */
            {8'h00}, /* 0xf1d7 */
            {8'h00}, /* 0xf1d6 */
            {8'h00}, /* 0xf1d5 */
            {8'h00}, /* 0xf1d4 */
            {8'h00}, /* 0xf1d3 */
            {8'h00}, /* 0xf1d2 */
            {8'h00}, /* 0xf1d1 */
            {8'h00}, /* 0xf1d0 */
            {8'h00}, /* 0xf1cf */
            {8'h00}, /* 0xf1ce */
            {8'h00}, /* 0xf1cd */
            {8'h00}, /* 0xf1cc */
            {8'h00}, /* 0xf1cb */
            {8'h00}, /* 0xf1ca */
            {8'h00}, /* 0xf1c9 */
            {8'h00}, /* 0xf1c8 */
            {8'h00}, /* 0xf1c7 */
            {8'h00}, /* 0xf1c6 */
            {8'h00}, /* 0xf1c5 */
            {8'h00}, /* 0xf1c4 */
            {8'h00}, /* 0xf1c3 */
            {8'h00}, /* 0xf1c2 */
            {8'h00}, /* 0xf1c1 */
            {8'h00}, /* 0xf1c0 */
            {8'h00}, /* 0xf1bf */
            {8'h00}, /* 0xf1be */
            {8'h00}, /* 0xf1bd */
            {8'h00}, /* 0xf1bc */
            {8'h00}, /* 0xf1bb */
            {8'h00}, /* 0xf1ba */
            {8'h00}, /* 0xf1b9 */
            {8'h00}, /* 0xf1b8 */
            {8'h00}, /* 0xf1b7 */
            {8'h00}, /* 0xf1b6 */
            {8'h00}, /* 0xf1b5 */
            {8'h00}, /* 0xf1b4 */
            {8'h00}, /* 0xf1b3 */
            {8'h00}, /* 0xf1b2 */
            {8'h00}, /* 0xf1b1 */
            {8'h00}, /* 0xf1b0 */
            {8'h00}, /* 0xf1af */
            {8'h00}, /* 0xf1ae */
            {8'h00}, /* 0xf1ad */
            {8'h00}, /* 0xf1ac */
            {8'h00}, /* 0xf1ab */
            {8'h00}, /* 0xf1aa */
            {8'h00}, /* 0xf1a9 */
            {8'h00}, /* 0xf1a8 */
            {8'h00}, /* 0xf1a7 */
            {8'h00}, /* 0xf1a6 */
            {8'h00}, /* 0xf1a5 */
            {8'h00}, /* 0xf1a4 */
            {8'h00}, /* 0xf1a3 */
            {8'h00}, /* 0xf1a2 */
            {8'h00}, /* 0xf1a1 */
            {8'h00}, /* 0xf1a0 */
            {8'h00}, /* 0xf19f */
            {8'h00}, /* 0xf19e */
            {8'h00}, /* 0xf19d */
            {8'h00}, /* 0xf19c */
            {8'h00}, /* 0xf19b */
            {8'h00}, /* 0xf19a */
            {8'h00}, /* 0xf199 */
            {8'h00}, /* 0xf198 */
            {8'h00}, /* 0xf197 */
            {8'h00}, /* 0xf196 */
            {8'h00}, /* 0xf195 */
            {8'h00}, /* 0xf194 */
            {8'h00}, /* 0xf193 */
            {8'h00}, /* 0xf192 */
            {8'h00}, /* 0xf191 */
            {8'h00}, /* 0xf190 */
            {8'h00}, /* 0xf18f */
            {8'h00}, /* 0xf18e */
            {8'h00}, /* 0xf18d */
            {8'h00}, /* 0xf18c */
            {8'h00}, /* 0xf18b */
            {8'h00}, /* 0xf18a */
            {8'h00}, /* 0xf189 */
            {8'h00}, /* 0xf188 */
            {8'h00}, /* 0xf187 */
            {8'h00}, /* 0xf186 */
            {8'h00}, /* 0xf185 */
            {8'h00}, /* 0xf184 */
            {8'h00}, /* 0xf183 */
            {8'h00}, /* 0xf182 */
            {8'h00}, /* 0xf181 */
            {8'h00}, /* 0xf180 */
            {8'h00}, /* 0xf17f */
            {8'h00}, /* 0xf17e */
            {8'h00}, /* 0xf17d */
            {8'h00}, /* 0xf17c */
            {8'h00}, /* 0xf17b */
            {8'h00}, /* 0xf17a */
            {8'h00}, /* 0xf179 */
            {8'h00}, /* 0xf178 */
            {8'h00}, /* 0xf177 */
            {8'h00}, /* 0xf176 */
            {8'h00}, /* 0xf175 */
            {8'h00}, /* 0xf174 */
            {8'h00}, /* 0xf173 */
            {8'h00}, /* 0xf172 */
            {8'h00}, /* 0xf171 */
            {8'h00}, /* 0xf170 */
            {8'h00}, /* 0xf16f */
            {8'h00}, /* 0xf16e */
            {8'h00}, /* 0xf16d */
            {8'h00}, /* 0xf16c */
            {8'h00}, /* 0xf16b */
            {8'h00}, /* 0xf16a */
            {8'h00}, /* 0xf169 */
            {8'h00}, /* 0xf168 */
            {8'h00}, /* 0xf167 */
            {8'h00}, /* 0xf166 */
            {8'h00}, /* 0xf165 */
            {8'h00}, /* 0xf164 */
            {8'h00}, /* 0xf163 */
            {8'h00}, /* 0xf162 */
            {8'h00}, /* 0xf161 */
            {8'h00}, /* 0xf160 */
            {8'h00}, /* 0xf15f */
            {8'h00}, /* 0xf15e */
            {8'h00}, /* 0xf15d */
            {8'h00}, /* 0xf15c */
            {8'h00}, /* 0xf15b */
            {8'h00}, /* 0xf15a */
            {8'h00}, /* 0xf159 */
            {8'h00}, /* 0xf158 */
            {8'h00}, /* 0xf157 */
            {8'h00}, /* 0xf156 */
            {8'h00}, /* 0xf155 */
            {8'h00}, /* 0xf154 */
            {8'h00}, /* 0xf153 */
            {8'h00}, /* 0xf152 */
            {8'h00}, /* 0xf151 */
            {8'h00}, /* 0xf150 */
            {8'h00}, /* 0xf14f */
            {8'h00}, /* 0xf14e */
            {8'h00}, /* 0xf14d */
            {8'h00}, /* 0xf14c */
            {8'h00}, /* 0xf14b */
            {8'h00}, /* 0xf14a */
            {8'h00}, /* 0xf149 */
            {8'h00}, /* 0xf148 */
            {8'h00}, /* 0xf147 */
            {8'h00}, /* 0xf146 */
            {8'h00}, /* 0xf145 */
            {8'h00}, /* 0xf144 */
            {8'h00}, /* 0xf143 */
            {8'h00}, /* 0xf142 */
            {8'h00}, /* 0xf141 */
            {8'h00}, /* 0xf140 */
            {8'h00}, /* 0xf13f */
            {8'h00}, /* 0xf13e */
            {8'h00}, /* 0xf13d */
            {8'h00}, /* 0xf13c */
            {8'h00}, /* 0xf13b */
            {8'h00}, /* 0xf13a */
            {8'h00}, /* 0xf139 */
            {8'h00}, /* 0xf138 */
            {8'h00}, /* 0xf137 */
            {8'h00}, /* 0xf136 */
            {8'h00}, /* 0xf135 */
            {8'h00}, /* 0xf134 */
            {8'h00}, /* 0xf133 */
            {8'h00}, /* 0xf132 */
            {8'h00}, /* 0xf131 */
            {8'h00}, /* 0xf130 */
            {8'h00}, /* 0xf12f */
            {8'h00}, /* 0xf12e */
            {8'h00}, /* 0xf12d */
            {8'h00}, /* 0xf12c */
            {8'h00}, /* 0xf12b */
            {8'h00}, /* 0xf12a */
            {8'h00}, /* 0xf129 */
            {8'h00}, /* 0xf128 */
            {8'h00}, /* 0xf127 */
            {8'h00}, /* 0xf126 */
            {8'h00}, /* 0xf125 */
            {8'h00}, /* 0xf124 */
            {8'h00}, /* 0xf123 */
            {8'h00}, /* 0xf122 */
            {8'h00}, /* 0xf121 */
            {8'h00}, /* 0xf120 */
            {8'h00}, /* 0xf11f */
            {8'h00}, /* 0xf11e */
            {8'h00}, /* 0xf11d */
            {8'h00}, /* 0xf11c */
            {8'h00}, /* 0xf11b */
            {8'h00}, /* 0xf11a */
            {8'h00}, /* 0xf119 */
            {8'h00}, /* 0xf118 */
            {8'h00}, /* 0xf117 */
            {8'h00}, /* 0xf116 */
            {8'h00}, /* 0xf115 */
            {8'h00}, /* 0xf114 */
            {8'h00}, /* 0xf113 */
            {8'h00}, /* 0xf112 */
            {8'h00}, /* 0xf111 */
            {8'h00}, /* 0xf110 */
            {8'h00}, /* 0xf10f */
            {8'h00}, /* 0xf10e */
            {8'h00}, /* 0xf10d */
            {8'h00}, /* 0xf10c */
            {8'h00}, /* 0xf10b */
            {8'h00}, /* 0xf10a */
            {8'h00}, /* 0xf109 */
            {8'h00}, /* 0xf108 */
            {8'h00}, /* 0xf107 */
            {8'h00}, /* 0xf106 */
            {8'h00}, /* 0xf105 */
            {8'h00}, /* 0xf104 */
            {8'h00}, /* 0xf103 */
            {8'h00}, /* 0xf102 */
            {8'h00}, /* 0xf101 */
            {8'h00}, /* 0xf100 */
            {8'h00}, /* 0xf0ff */
            {8'h00}, /* 0xf0fe */
            {8'h00}, /* 0xf0fd */
            {8'h00}, /* 0xf0fc */
            {8'h00}, /* 0xf0fb */
            {8'h00}, /* 0xf0fa */
            {8'h00}, /* 0xf0f9 */
            {8'h00}, /* 0xf0f8 */
            {8'h00}, /* 0xf0f7 */
            {8'h00}, /* 0xf0f6 */
            {8'h00}, /* 0xf0f5 */
            {8'h00}, /* 0xf0f4 */
            {8'h00}, /* 0xf0f3 */
            {8'h00}, /* 0xf0f2 */
            {8'h00}, /* 0xf0f1 */
            {8'h00}, /* 0xf0f0 */
            {8'h00}, /* 0xf0ef */
            {8'h00}, /* 0xf0ee */
            {8'h00}, /* 0xf0ed */
            {8'h00}, /* 0xf0ec */
            {8'h00}, /* 0xf0eb */
            {8'h00}, /* 0xf0ea */
            {8'h00}, /* 0xf0e9 */
            {8'h00}, /* 0xf0e8 */
            {8'h00}, /* 0xf0e7 */
            {8'h00}, /* 0xf0e6 */
            {8'h00}, /* 0xf0e5 */
            {8'h00}, /* 0xf0e4 */
            {8'h00}, /* 0xf0e3 */
            {8'h00}, /* 0xf0e2 */
            {8'h00}, /* 0xf0e1 */
            {8'h00}, /* 0xf0e0 */
            {8'h00}, /* 0xf0df */
            {8'h00}, /* 0xf0de */
            {8'h00}, /* 0xf0dd */
            {8'h00}, /* 0xf0dc */
            {8'h00}, /* 0xf0db */
            {8'h00}, /* 0xf0da */
            {8'h00}, /* 0xf0d9 */
            {8'h00}, /* 0xf0d8 */
            {8'h00}, /* 0xf0d7 */
            {8'h00}, /* 0xf0d6 */
            {8'h00}, /* 0xf0d5 */
            {8'h00}, /* 0xf0d4 */
            {8'h00}, /* 0xf0d3 */
            {8'h00}, /* 0xf0d2 */
            {8'h00}, /* 0xf0d1 */
            {8'h00}, /* 0xf0d0 */
            {8'h00}, /* 0xf0cf */
            {8'h00}, /* 0xf0ce */
            {8'h00}, /* 0xf0cd */
            {8'h00}, /* 0xf0cc */
            {8'h00}, /* 0xf0cb */
            {8'h00}, /* 0xf0ca */
            {8'h00}, /* 0xf0c9 */
            {8'h00}, /* 0xf0c8 */
            {8'h00}, /* 0xf0c7 */
            {8'h00}, /* 0xf0c6 */
            {8'h00}, /* 0xf0c5 */
            {8'h00}, /* 0xf0c4 */
            {8'h00}, /* 0xf0c3 */
            {8'h00}, /* 0xf0c2 */
            {8'h00}, /* 0xf0c1 */
            {8'h00}, /* 0xf0c0 */
            {8'h00}, /* 0xf0bf */
            {8'h00}, /* 0xf0be */
            {8'h00}, /* 0xf0bd */
            {8'h00}, /* 0xf0bc */
            {8'h00}, /* 0xf0bb */
            {8'h00}, /* 0xf0ba */
            {8'h00}, /* 0xf0b9 */
            {8'h00}, /* 0xf0b8 */
            {8'h00}, /* 0xf0b7 */
            {8'h00}, /* 0xf0b6 */
            {8'h00}, /* 0xf0b5 */
            {8'h00}, /* 0xf0b4 */
            {8'h00}, /* 0xf0b3 */
            {8'h00}, /* 0xf0b2 */
            {8'h00}, /* 0xf0b1 */
            {8'h00}, /* 0xf0b0 */
            {8'h00}, /* 0xf0af */
            {8'h00}, /* 0xf0ae */
            {8'h00}, /* 0xf0ad */
            {8'h00}, /* 0xf0ac */
            {8'h00}, /* 0xf0ab */
            {8'h00}, /* 0xf0aa */
            {8'h00}, /* 0xf0a9 */
            {8'h00}, /* 0xf0a8 */
            {8'h00}, /* 0xf0a7 */
            {8'h00}, /* 0xf0a6 */
            {8'h00}, /* 0xf0a5 */
            {8'h00}, /* 0xf0a4 */
            {8'h00}, /* 0xf0a3 */
            {8'h00}, /* 0xf0a2 */
            {8'h00}, /* 0xf0a1 */
            {8'h00}, /* 0xf0a0 */
            {8'h00}, /* 0xf09f */
            {8'h00}, /* 0xf09e */
            {8'h00}, /* 0xf09d */
            {8'h00}, /* 0xf09c */
            {8'h00}, /* 0xf09b */
            {8'h00}, /* 0xf09a */
            {8'h00}, /* 0xf099 */
            {8'h00}, /* 0xf098 */
            {8'h00}, /* 0xf097 */
            {8'h00}, /* 0xf096 */
            {8'h00}, /* 0xf095 */
            {8'h00}, /* 0xf094 */
            {8'h00}, /* 0xf093 */
            {8'h00}, /* 0xf092 */
            {8'h00}, /* 0xf091 */
            {8'h00}, /* 0xf090 */
            {8'h00}, /* 0xf08f */
            {8'h00}, /* 0xf08e */
            {8'h00}, /* 0xf08d */
            {8'h00}, /* 0xf08c */
            {8'h00}, /* 0xf08b */
            {8'h00}, /* 0xf08a */
            {8'h00}, /* 0xf089 */
            {8'h00}, /* 0xf088 */
            {8'h00}, /* 0xf087 */
            {8'h00}, /* 0xf086 */
            {8'h00}, /* 0xf085 */
            {8'h00}, /* 0xf084 */
            {8'h00}, /* 0xf083 */
            {8'h00}, /* 0xf082 */
            {8'h00}, /* 0xf081 */
            {8'h00}, /* 0xf080 */
            {8'h00}, /* 0xf07f */
            {8'h00}, /* 0xf07e */
            {8'h00}, /* 0xf07d */
            {8'h00}, /* 0xf07c */
            {8'h00}, /* 0xf07b */
            {8'h00}, /* 0xf07a */
            {8'h00}, /* 0xf079 */
            {8'h00}, /* 0xf078 */
            {8'h00}, /* 0xf077 */
            {8'h00}, /* 0xf076 */
            {8'h00}, /* 0xf075 */
            {8'h00}, /* 0xf074 */
            {8'h00}, /* 0xf073 */
            {8'h00}, /* 0xf072 */
            {8'h00}, /* 0xf071 */
            {8'h00}, /* 0xf070 */
            {8'h00}, /* 0xf06f */
            {8'h00}, /* 0xf06e */
            {8'h00}, /* 0xf06d */
            {8'h00}, /* 0xf06c */
            {8'h00}, /* 0xf06b */
            {8'h00}, /* 0xf06a */
            {8'h00}, /* 0xf069 */
            {8'h00}, /* 0xf068 */
            {8'h00}, /* 0xf067 */
            {8'h00}, /* 0xf066 */
            {8'h00}, /* 0xf065 */
            {8'h00}, /* 0xf064 */
            {8'h00}, /* 0xf063 */
            {8'h00}, /* 0xf062 */
            {8'h00}, /* 0xf061 */
            {8'h00}, /* 0xf060 */
            {8'h00}, /* 0xf05f */
            {8'h00}, /* 0xf05e */
            {8'h00}, /* 0xf05d */
            {8'h00}, /* 0xf05c */
            {8'h00}, /* 0xf05b */
            {8'h00}, /* 0xf05a */
            {8'h00}, /* 0xf059 */
            {8'h00}, /* 0xf058 */
            {8'h00}, /* 0xf057 */
            {8'h00}, /* 0xf056 */
            {8'h00}, /* 0xf055 */
            {8'h00}, /* 0xf054 */
            {8'h00}, /* 0xf053 */
            {8'h00}, /* 0xf052 */
            {8'h00}, /* 0xf051 */
            {8'h00}, /* 0xf050 */
            {8'h00}, /* 0xf04f */
            {8'h00}, /* 0xf04e */
            {8'h00}, /* 0xf04d */
            {8'h00}, /* 0xf04c */
            {8'h00}, /* 0xf04b */
            {8'h00}, /* 0xf04a */
            {8'h00}, /* 0xf049 */
            {8'h00}, /* 0xf048 */
            {8'h00}, /* 0xf047 */
            {8'h00}, /* 0xf046 */
            {8'h00}, /* 0xf045 */
            {8'h00}, /* 0xf044 */
            {8'h00}, /* 0xf043 */
            {8'h00}, /* 0xf042 */
            {8'h00}, /* 0xf041 */
            {8'h00}, /* 0xf040 */
            {8'h00}, /* 0xf03f */
            {8'h00}, /* 0xf03e */
            {8'h00}, /* 0xf03d */
            {8'h00}, /* 0xf03c */
            {8'h00}, /* 0xf03b */
            {8'h00}, /* 0xf03a */
            {8'h00}, /* 0xf039 */
            {8'h00}, /* 0xf038 */
            {8'h00}, /* 0xf037 */
            {8'h00}, /* 0xf036 */
            {8'h00}, /* 0xf035 */
            {8'h00}, /* 0xf034 */
            {8'h00}, /* 0xf033 */
            {8'h00}, /* 0xf032 */
            {8'h00}, /* 0xf031 */
            {8'h00}, /* 0xf030 */
            {8'h00}, /* 0xf02f */
            {8'h00}, /* 0xf02e */
            {8'h00}, /* 0xf02d */
            {8'h00}, /* 0xf02c */
            {8'h00}, /* 0xf02b */
            {8'h00}, /* 0xf02a */
            {8'h00}, /* 0xf029 */
            {8'h00}, /* 0xf028 */
            {8'h00}, /* 0xf027 */
            {8'h00}, /* 0xf026 */
            {8'h00}, /* 0xf025 */
            {8'h00}, /* 0xf024 */
            {8'h00}, /* 0xf023 */
            {8'h00}, /* 0xf022 */
            {8'h00}, /* 0xf021 */
            {8'h00}, /* 0xf020 */
            {8'h00}, /* 0xf01f */
            {8'h00}, /* 0xf01e */
            {8'h00}, /* 0xf01d */
            {8'h00}, /* 0xf01c */
            {8'h00}, /* 0xf01b */
            {8'h00}, /* 0xf01a */
            {8'h00}, /* 0xf019 */
            {8'h00}, /* 0xf018 */
            {8'h00}, /* 0xf017 */
            {8'h00}, /* 0xf016 */
            {8'h00}, /* 0xf015 */
            {8'h00}, /* 0xf014 */
            {8'h00}, /* 0xf013 */
            {8'h00}, /* 0xf012 */
            {8'h00}, /* 0xf011 */
            {8'h00}, /* 0xf010 */
            {8'h00}, /* 0xf00f */
            {8'h00}, /* 0xf00e */
            {8'h00}, /* 0xf00d */
            {8'h00}, /* 0xf00c */
            {8'h00}, /* 0xf00b */
            {8'h00}, /* 0xf00a */
            {8'h00}, /* 0xf009 */
            {8'h00}, /* 0xf008 */
            {8'h00}, /* 0xf007 */
            {8'h00}, /* 0xf006 */
            {8'h00}, /* 0xf005 */
            {8'h00}, /* 0xf004 */
            {8'h00}, /* 0xf003 */
            {8'h00}, /* 0xf002 */
            {8'h00}, /* 0xf001 */
            {8'h00}, /* 0xf000 */
            {8'h00}, /* 0xefff */
            {8'h00}, /* 0xeffe */
            {8'h00}, /* 0xeffd */
            {8'h00}, /* 0xeffc */
            {8'h00}, /* 0xeffb */
            {8'h00}, /* 0xeffa */
            {8'h00}, /* 0xeff9 */
            {8'h00}, /* 0xeff8 */
            {8'h00}, /* 0xeff7 */
            {8'h00}, /* 0xeff6 */
            {8'h00}, /* 0xeff5 */
            {8'h00}, /* 0xeff4 */
            {8'h00}, /* 0xeff3 */
            {8'h00}, /* 0xeff2 */
            {8'h00}, /* 0xeff1 */
            {8'h00}, /* 0xeff0 */
            {8'h00}, /* 0xefef */
            {8'h00}, /* 0xefee */
            {8'h00}, /* 0xefed */
            {8'h00}, /* 0xefec */
            {8'h00}, /* 0xefeb */
            {8'h00}, /* 0xefea */
            {8'h00}, /* 0xefe9 */
            {8'h00}, /* 0xefe8 */
            {8'h00}, /* 0xefe7 */
            {8'h00}, /* 0xefe6 */
            {8'h00}, /* 0xefe5 */
            {8'h00}, /* 0xefe4 */
            {8'h00}, /* 0xefe3 */
            {8'h00}, /* 0xefe2 */
            {8'h00}, /* 0xefe1 */
            {8'h00}, /* 0xefe0 */
            {8'h00}, /* 0xefdf */
            {8'h00}, /* 0xefde */
            {8'h00}, /* 0xefdd */
            {8'h00}, /* 0xefdc */
            {8'h00}, /* 0xefdb */
            {8'h00}, /* 0xefda */
            {8'h00}, /* 0xefd9 */
            {8'h00}, /* 0xefd8 */
            {8'h00}, /* 0xefd7 */
            {8'h00}, /* 0xefd6 */
            {8'h00}, /* 0xefd5 */
            {8'h00}, /* 0xefd4 */
            {8'h00}, /* 0xefd3 */
            {8'h00}, /* 0xefd2 */
            {8'h00}, /* 0xefd1 */
            {8'h00}, /* 0xefd0 */
            {8'h00}, /* 0xefcf */
            {8'h00}, /* 0xefce */
            {8'h00}, /* 0xefcd */
            {8'h00}, /* 0xefcc */
            {8'h00}, /* 0xefcb */
            {8'h00}, /* 0xefca */
            {8'h00}, /* 0xefc9 */
            {8'h00}, /* 0xefc8 */
            {8'h00}, /* 0xefc7 */
            {8'h00}, /* 0xefc6 */
            {8'h00}, /* 0xefc5 */
            {8'h00}, /* 0xefc4 */
            {8'h00}, /* 0xefc3 */
            {8'h00}, /* 0xefc2 */
            {8'h00}, /* 0xefc1 */
            {8'h00}, /* 0xefc0 */
            {8'h00}, /* 0xefbf */
            {8'h00}, /* 0xefbe */
            {8'h00}, /* 0xefbd */
            {8'h00}, /* 0xefbc */
            {8'h00}, /* 0xefbb */
            {8'h00}, /* 0xefba */
            {8'h00}, /* 0xefb9 */
            {8'h00}, /* 0xefb8 */
            {8'h00}, /* 0xefb7 */
            {8'h00}, /* 0xefb6 */
            {8'h00}, /* 0xefb5 */
            {8'h00}, /* 0xefb4 */
            {8'h00}, /* 0xefb3 */
            {8'h00}, /* 0xefb2 */
            {8'h00}, /* 0xefb1 */
            {8'h00}, /* 0xefb0 */
            {8'h00}, /* 0xefaf */
            {8'h00}, /* 0xefae */
            {8'h00}, /* 0xefad */
            {8'h00}, /* 0xefac */
            {8'h00}, /* 0xefab */
            {8'h00}, /* 0xefaa */
            {8'h00}, /* 0xefa9 */
            {8'h00}, /* 0xefa8 */
            {8'h00}, /* 0xefa7 */
            {8'h00}, /* 0xefa6 */
            {8'h00}, /* 0xefa5 */
            {8'h00}, /* 0xefa4 */
            {8'h00}, /* 0xefa3 */
            {8'h00}, /* 0xefa2 */
            {8'h00}, /* 0xefa1 */
            {8'h00}, /* 0xefa0 */
            {8'h00}, /* 0xef9f */
            {8'h00}, /* 0xef9e */
            {8'h00}, /* 0xef9d */
            {8'h00}, /* 0xef9c */
            {8'h00}, /* 0xef9b */
            {8'h00}, /* 0xef9a */
            {8'h00}, /* 0xef99 */
            {8'h00}, /* 0xef98 */
            {8'h00}, /* 0xef97 */
            {8'h00}, /* 0xef96 */
            {8'h00}, /* 0xef95 */
            {8'h00}, /* 0xef94 */
            {8'h00}, /* 0xef93 */
            {8'h00}, /* 0xef92 */
            {8'h00}, /* 0xef91 */
            {8'h00}, /* 0xef90 */
            {8'h00}, /* 0xef8f */
            {8'h00}, /* 0xef8e */
            {8'h00}, /* 0xef8d */
            {8'h00}, /* 0xef8c */
            {8'h00}, /* 0xef8b */
            {8'h00}, /* 0xef8a */
            {8'h00}, /* 0xef89 */
            {8'h00}, /* 0xef88 */
            {8'h00}, /* 0xef87 */
            {8'h00}, /* 0xef86 */
            {8'h00}, /* 0xef85 */
            {8'h00}, /* 0xef84 */
            {8'h00}, /* 0xef83 */
            {8'h00}, /* 0xef82 */
            {8'h00}, /* 0xef81 */
            {8'h00}, /* 0xef80 */
            {8'h00}, /* 0xef7f */
            {8'h00}, /* 0xef7e */
            {8'h00}, /* 0xef7d */
            {8'h00}, /* 0xef7c */
            {8'h00}, /* 0xef7b */
            {8'h00}, /* 0xef7a */
            {8'h00}, /* 0xef79 */
            {8'h00}, /* 0xef78 */
            {8'h00}, /* 0xef77 */
            {8'h00}, /* 0xef76 */
            {8'h00}, /* 0xef75 */
            {8'h00}, /* 0xef74 */
            {8'h00}, /* 0xef73 */
            {8'h00}, /* 0xef72 */
            {8'h00}, /* 0xef71 */
            {8'h00}, /* 0xef70 */
            {8'h00}, /* 0xef6f */
            {8'h00}, /* 0xef6e */
            {8'h00}, /* 0xef6d */
            {8'h00}, /* 0xef6c */
            {8'h00}, /* 0xef6b */
            {8'h00}, /* 0xef6a */
            {8'h00}, /* 0xef69 */
            {8'h00}, /* 0xef68 */
            {8'h00}, /* 0xef67 */
            {8'h00}, /* 0xef66 */
            {8'h00}, /* 0xef65 */
            {8'h00}, /* 0xef64 */
            {8'h00}, /* 0xef63 */
            {8'h00}, /* 0xef62 */
            {8'h00}, /* 0xef61 */
            {8'h00}, /* 0xef60 */
            {8'h00}, /* 0xef5f */
            {8'h00}, /* 0xef5e */
            {8'h00}, /* 0xef5d */
            {8'h00}, /* 0xef5c */
            {8'h00}, /* 0xef5b */
            {8'h00}, /* 0xef5a */
            {8'h00}, /* 0xef59 */
            {8'h00}, /* 0xef58 */
            {8'h00}, /* 0xef57 */
            {8'h00}, /* 0xef56 */
            {8'h00}, /* 0xef55 */
            {8'h00}, /* 0xef54 */
            {8'h00}, /* 0xef53 */
            {8'h00}, /* 0xef52 */
            {8'h00}, /* 0xef51 */
            {8'h00}, /* 0xef50 */
            {8'h00}, /* 0xef4f */
            {8'h00}, /* 0xef4e */
            {8'h00}, /* 0xef4d */
            {8'h00}, /* 0xef4c */
            {8'h00}, /* 0xef4b */
            {8'h00}, /* 0xef4a */
            {8'h00}, /* 0xef49 */
            {8'h00}, /* 0xef48 */
            {8'h00}, /* 0xef47 */
            {8'h00}, /* 0xef46 */
            {8'h00}, /* 0xef45 */
            {8'h00}, /* 0xef44 */
            {8'h00}, /* 0xef43 */
            {8'h00}, /* 0xef42 */
            {8'h00}, /* 0xef41 */
            {8'h00}, /* 0xef40 */
            {8'h00}, /* 0xef3f */
            {8'h00}, /* 0xef3e */
            {8'h00}, /* 0xef3d */
            {8'h00}, /* 0xef3c */
            {8'h00}, /* 0xef3b */
            {8'h00}, /* 0xef3a */
            {8'h00}, /* 0xef39 */
            {8'h00}, /* 0xef38 */
            {8'h00}, /* 0xef37 */
            {8'h00}, /* 0xef36 */
            {8'h00}, /* 0xef35 */
            {8'h00}, /* 0xef34 */
            {8'h00}, /* 0xef33 */
            {8'h00}, /* 0xef32 */
            {8'h00}, /* 0xef31 */
            {8'h00}, /* 0xef30 */
            {8'h00}, /* 0xef2f */
            {8'h00}, /* 0xef2e */
            {8'h00}, /* 0xef2d */
            {8'h00}, /* 0xef2c */
            {8'h00}, /* 0xef2b */
            {8'h00}, /* 0xef2a */
            {8'h00}, /* 0xef29 */
            {8'h00}, /* 0xef28 */
            {8'h00}, /* 0xef27 */
            {8'h00}, /* 0xef26 */
            {8'h00}, /* 0xef25 */
            {8'h00}, /* 0xef24 */
            {8'h00}, /* 0xef23 */
            {8'h00}, /* 0xef22 */
            {8'h00}, /* 0xef21 */
            {8'h00}, /* 0xef20 */
            {8'h00}, /* 0xef1f */
            {8'h00}, /* 0xef1e */
            {8'h00}, /* 0xef1d */
            {8'h00}, /* 0xef1c */
            {8'h00}, /* 0xef1b */
            {8'h00}, /* 0xef1a */
            {8'h00}, /* 0xef19 */
            {8'h00}, /* 0xef18 */
            {8'h00}, /* 0xef17 */
            {8'h00}, /* 0xef16 */
            {8'h00}, /* 0xef15 */
            {8'h00}, /* 0xef14 */
            {8'h00}, /* 0xef13 */
            {8'h00}, /* 0xef12 */
            {8'h00}, /* 0xef11 */
            {8'h00}, /* 0xef10 */
            {8'h00}, /* 0xef0f */
            {8'h00}, /* 0xef0e */
            {8'h00}, /* 0xef0d */
            {8'h00}, /* 0xef0c */
            {8'h00}, /* 0xef0b */
            {8'h00}, /* 0xef0a */
            {8'h00}, /* 0xef09 */
            {8'h00}, /* 0xef08 */
            {8'h00}, /* 0xef07 */
            {8'h00}, /* 0xef06 */
            {8'h00}, /* 0xef05 */
            {8'h00}, /* 0xef04 */
            {8'h00}, /* 0xef03 */
            {8'h00}, /* 0xef02 */
            {8'h00}, /* 0xef01 */
            {8'h00}, /* 0xef00 */
            {8'h00}, /* 0xeeff */
            {8'h00}, /* 0xeefe */
            {8'h00}, /* 0xeefd */
            {8'h00}, /* 0xeefc */
            {8'h00}, /* 0xeefb */
            {8'h00}, /* 0xeefa */
            {8'h00}, /* 0xeef9 */
            {8'h00}, /* 0xeef8 */
            {8'h00}, /* 0xeef7 */
            {8'h00}, /* 0xeef6 */
            {8'h00}, /* 0xeef5 */
            {8'h00}, /* 0xeef4 */
            {8'h00}, /* 0xeef3 */
            {8'h00}, /* 0xeef2 */
            {8'h00}, /* 0xeef1 */
            {8'h00}, /* 0xeef0 */
            {8'h00}, /* 0xeeef */
            {8'h00}, /* 0xeeee */
            {8'h00}, /* 0xeeed */
            {8'h00}, /* 0xeeec */
            {8'h00}, /* 0xeeeb */
            {8'h00}, /* 0xeeea */
            {8'h00}, /* 0xeee9 */
            {8'h00}, /* 0xeee8 */
            {8'h00}, /* 0xeee7 */
            {8'h00}, /* 0xeee6 */
            {8'h00}, /* 0xeee5 */
            {8'h00}, /* 0xeee4 */
            {8'h00}, /* 0xeee3 */
            {8'h00}, /* 0xeee2 */
            {8'h00}, /* 0xeee1 */
            {8'h00}, /* 0xeee0 */
            {8'h00}, /* 0xeedf */
            {8'h00}, /* 0xeede */
            {8'h00}, /* 0xeedd */
            {8'h00}, /* 0xeedc */
            {8'h00}, /* 0xeedb */
            {8'h00}, /* 0xeeda */
            {8'h00}, /* 0xeed9 */
            {8'h00}, /* 0xeed8 */
            {8'h00}, /* 0xeed7 */
            {8'h00}, /* 0xeed6 */
            {8'h00}, /* 0xeed5 */
            {8'h00}, /* 0xeed4 */
            {8'h00}, /* 0xeed3 */
            {8'h00}, /* 0xeed2 */
            {8'h00}, /* 0xeed1 */
            {8'h00}, /* 0xeed0 */
            {8'h00}, /* 0xeecf */
            {8'h00}, /* 0xeece */
            {8'h00}, /* 0xeecd */
            {8'h00}, /* 0xeecc */
            {8'h00}, /* 0xeecb */
            {8'h00}, /* 0xeeca */
            {8'h00}, /* 0xeec9 */
            {8'h00}, /* 0xeec8 */
            {8'h00}, /* 0xeec7 */
            {8'h00}, /* 0xeec6 */
            {8'h00}, /* 0xeec5 */
            {8'h00}, /* 0xeec4 */
            {8'h00}, /* 0xeec3 */
            {8'h00}, /* 0xeec2 */
            {8'h00}, /* 0xeec1 */
            {8'h00}, /* 0xeec0 */
            {8'h00}, /* 0xeebf */
            {8'h00}, /* 0xeebe */
            {8'h00}, /* 0xeebd */
            {8'h00}, /* 0xeebc */
            {8'h00}, /* 0xeebb */
            {8'h00}, /* 0xeeba */
            {8'h00}, /* 0xeeb9 */
            {8'h00}, /* 0xeeb8 */
            {8'h00}, /* 0xeeb7 */
            {8'h00}, /* 0xeeb6 */
            {8'h00}, /* 0xeeb5 */
            {8'h00}, /* 0xeeb4 */
            {8'h00}, /* 0xeeb3 */
            {8'h00}, /* 0xeeb2 */
            {8'h00}, /* 0xeeb1 */
            {8'h00}, /* 0xeeb0 */
            {8'h00}, /* 0xeeaf */
            {8'h00}, /* 0xeeae */
            {8'h00}, /* 0xeead */
            {8'h00}, /* 0xeeac */
            {8'h00}, /* 0xeeab */
            {8'h00}, /* 0xeeaa */
            {8'h00}, /* 0xeea9 */
            {8'h00}, /* 0xeea8 */
            {8'h00}, /* 0xeea7 */
            {8'h00}, /* 0xeea6 */
            {8'h00}, /* 0xeea5 */
            {8'h00}, /* 0xeea4 */
            {8'h00}, /* 0xeea3 */
            {8'h00}, /* 0xeea2 */
            {8'h00}, /* 0xeea1 */
            {8'h00}, /* 0xeea0 */
            {8'h00}, /* 0xee9f */
            {8'h00}, /* 0xee9e */
            {8'h00}, /* 0xee9d */
            {8'h00}, /* 0xee9c */
            {8'h00}, /* 0xee9b */
            {8'h00}, /* 0xee9a */
            {8'h00}, /* 0xee99 */
            {8'h00}, /* 0xee98 */
            {8'h00}, /* 0xee97 */
            {8'h00}, /* 0xee96 */
            {8'h00}, /* 0xee95 */
            {8'h00}, /* 0xee94 */
            {8'h00}, /* 0xee93 */
            {8'h00}, /* 0xee92 */
            {8'h00}, /* 0xee91 */
            {8'h00}, /* 0xee90 */
            {8'h00}, /* 0xee8f */
            {8'h00}, /* 0xee8e */
            {8'h00}, /* 0xee8d */
            {8'h00}, /* 0xee8c */
            {8'h00}, /* 0xee8b */
            {8'h00}, /* 0xee8a */
            {8'h00}, /* 0xee89 */
            {8'h00}, /* 0xee88 */
            {8'h00}, /* 0xee87 */
            {8'h00}, /* 0xee86 */
            {8'h00}, /* 0xee85 */
            {8'h00}, /* 0xee84 */
            {8'h00}, /* 0xee83 */
            {8'h00}, /* 0xee82 */
            {8'h00}, /* 0xee81 */
            {8'h00}, /* 0xee80 */
            {8'h00}, /* 0xee7f */
            {8'h00}, /* 0xee7e */
            {8'h00}, /* 0xee7d */
            {8'h00}, /* 0xee7c */
            {8'h00}, /* 0xee7b */
            {8'h00}, /* 0xee7a */
            {8'h00}, /* 0xee79 */
            {8'h00}, /* 0xee78 */
            {8'h00}, /* 0xee77 */
            {8'h00}, /* 0xee76 */
            {8'h00}, /* 0xee75 */
            {8'h00}, /* 0xee74 */
            {8'h00}, /* 0xee73 */
            {8'h00}, /* 0xee72 */
            {8'h00}, /* 0xee71 */
            {8'h00}, /* 0xee70 */
            {8'h00}, /* 0xee6f */
            {8'h00}, /* 0xee6e */
            {8'h00}, /* 0xee6d */
            {8'h00}, /* 0xee6c */
            {8'h00}, /* 0xee6b */
            {8'h00}, /* 0xee6a */
            {8'h00}, /* 0xee69 */
            {8'h00}, /* 0xee68 */
            {8'h00}, /* 0xee67 */
            {8'h00}, /* 0xee66 */
            {8'h00}, /* 0xee65 */
            {8'h00}, /* 0xee64 */
            {8'h00}, /* 0xee63 */
            {8'h00}, /* 0xee62 */
            {8'h00}, /* 0xee61 */
            {8'h00}, /* 0xee60 */
            {8'h00}, /* 0xee5f */
            {8'h00}, /* 0xee5e */
            {8'h00}, /* 0xee5d */
            {8'h00}, /* 0xee5c */
            {8'h00}, /* 0xee5b */
            {8'h00}, /* 0xee5a */
            {8'h00}, /* 0xee59 */
            {8'h00}, /* 0xee58 */
            {8'h00}, /* 0xee57 */
            {8'h00}, /* 0xee56 */
            {8'h00}, /* 0xee55 */
            {8'h00}, /* 0xee54 */
            {8'h00}, /* 0xee53 */
            {8'h00}, /* 0xee52 */
            {8'h00}, /* 0xee51 */
            {8'h00}, /* 0xee50 */
            {8'h00}, /* 0xee4f */
            {8'h00}, /* 0xee4e */
            {8'h00}, /* 0xee4d */
            {8'h00}, /* 0xee4c */
            {8'h00}, /* 0xee4b */
            {8'h00}, /* 0xee4a */
            {8'h00}, /* 0xee49 */
            {8'h00}, /* 0xee48 */
            {8'h00}, /* 0xee47 */
            {8'h00}, /* 0xee46 */
            {8'h00}, /* 0xee45 */
            {8'h00}, /* 0xee44 */
            {8'h00}, /* 0xee43 */
            {8'h00}, /* 0xee42 */
            {8'h00}, /* 0xee41 */
            {8'h00}, /* 0xee40 */
            {8'h00}, /* 0xee3f */
            {8'h00}, /* 0xee3e */
            {8'h00}, /* 0xee3d */
            {8'h00}, /* 0xee3c */
            {8'h00}, /* 0xee3b */
            {8'h00}, /* 0xee3a */
            {8'h00}, /* 0xee39 */
            {8'h00}, /* 0xee38 */
            {8'h00}, /* 0xee37 */
            {8'h00}, /* 0xee36 */
            {8'h00}, /* 0xee35 */
            {8'h00}, /* 0xee34 */
            {8'h00}, /* 0xee33 */
            {8'h00}, /* 0xee32 */
            {8'h00}, /* 0xee31 */
            {8'h00}, /* 0xee30 */
            {8'h00}, /* 0xee2f */
            {8'h00}, /* 0xee2e */
            {8'h00}, /* 0xee2d */
            {8'h00}, /* 0xee2c */
            {8'h00}, /* 0xee2b */
            {8'h00}, /* 0xee2a */
            {8'h00}, /* 0xee29 */
            {8'h00}, /* 0xee28 */
            {8'h00}, /* 0xee27 */
            {8'h00}, /* 0xee26 */
            {8'h00}, /* 0xee25 */
            {8'h00}, /* 0xee24 */
            {8'h00}, /* 0xee23 */
            {8'h00}, /* 0xee22 */
            {8'h00}, /* 0xee21 */
            {8'h00}, /* 0xee20 */
            {8'h00}, /* 0xee1f */
            {8'h00}, /* 0xee1e */
            {8'h00}, /* 0xee1d */
            {8'h00}, /* 0xee1c */
            {8'h00}, /* 0xee1b */
            {8'h00}, /* 0xee1a */
            {8'h00}, /* 0xee19 */
            {8'h00}, /* 0xee18 */
            {8'h00}, /* 0xee17 */
            {8'h00}, /* 0xee16 */
            {8'h00}, /* 0xee15 */
            {8'h00}, /* 0xee14 */
            {8'h00}, /* 0xee13 */
            {8'h00}, /* 0xee12 */
            {8'h00}, /* 0xee11 */
            {8'h00}, /* 0xee10 */
            {8'h00}, /* 0xee0f */
            {8'h00}, /* 0xee0e */
            {8'h00}, /* 0xee0d */
            {8'h00}, /* 0xee0c */
            {8'h00}, /* 0xee0b */
            {8'h00}, /* 0xee0a */
            {8'h00}, /* 0xee09 */
            {8'h00}, /* 0xee08 */
            {8'h00}, /* 0xee07 */
            {8'h00}, /* 0xee06 */
            {8'h00}, /* 0xee05 */
            {8'h00}, /* 0xee04 */
            {8'h00}, /* 0xee03 */
            {8'h00}, /* 0xee02 */
            {8'h00}, /* 0xee01 */
            {8'h00}, /* 0xee00 */
            {8'h00}, /* 0xedff */
            {8'h00}, /* 0xedfe */
            {8'h00}, /* 0xedfd */
            {8'h00}, /* 0xedfc */
            {8'h00}, /* 0xedfb */
            {8'h00}, /* 0xedfa */
            {8'h00}, /* 0xedf9 */
            {8'h00}, /* 0xedf8 */
            {8'h00}, /* 0xedf7 */
            {8'h00}, /* 0xedf6 */
            {8'h00}, /* 0xedf5 */
            {8'h00}, /* 0xedf4 */
            {8'h00}, /* 0xedf3 */
            {8'h00}, /* 0xedf2 */
            {8'h00}, /* 0xedf1 */
            {8'h00}, /* 0xedf0 */
            {8'h00}, /* 0xedef */
            {8'h00}, /* 0xedee */
            {8'h00}, /* 0xeded */
            {8'h00}, /* 0xedec */
            {8'h00}, /* 0xedeb */
            {8'h00}, /* 0xedea */
            {8'h00}, /* 0xede9 */
            {8'h00}, /* 0xede8 */
            {8'h00}, /* 0xede7 */
            {8'h00}, /* 0xede6 */
            {8'h00}, /* 0xede5 */
            {8'h00}, /* 0xede4 */
            {8'h00}, /* 0xede3 */
            {8'h00}, /* 0xede2 */
            {8'h00}, /* 0xede1 */
            {8'h00}, /* 0xede0 */
            {8'h00}, /* 0xeddf */
            {8'h00}, /* 0xedde */
            {8'h00}, /* 0xeddd */
            {8'h00}, /* 0xeddc */
            {8'h00}, /* 0xeddb */
            {8'h00}, /* 0xedda */
            {8'h00}, /* 0xedd9 */
            {8'h00}, /* 0xedd8 */
            {8'h00}, /* 0xedd7 */
            {8'h00}, /* 0xedd6 */
            {8'h00}, /* 0xedd5 */
            {8'h00}, /* 0xedd4 */
            {8'h00}, /* 0xedd3 */
            {8'h00}, /* 0xedd2 */
            {8'h00}, /* 0xedd1 */
            {8'h00}, /* 0xedd0 */
            {8'h00}, /* 0xedcf */
            {8'h00}, /* 0xedce */
            {8'h00}, /* 0xedcd */
            {8'h00}, /* 0xedcc */
            {8'h00}, /* 0xedcb */
            {8'h00}, /* 0xedca */
            {8'h00}, /* 0xedc9 */
            {8'h00}, /* 0xedc8 */
            {8'h00}, /* 0xedc7 */
            {8'h00}, /* 0xedc6 */
            {8'h00}, /* 0xedc5 */
            {8'h00}, /* 0xedc4 */
            {8'h00}, /* 0xedc3 */
            {8'h00}, /* 0xedc2 */
            {8'h00}, /* 0xedc1 */
            {8'h00}, /* 0xedc0 */
            {8'h00}, /* 0xedbf */
            {8'h00}, /* 0xedbe */
            {8'h00}, /* 0xedbd */
            {8'h00}, /* 0xedbc */
            {8'h00}, /* 0xedbb */
            {8'h00}, /* 0xedba */
            {8'h00}, /* 0xedb9 */
            {8'h00}, /* 0xedb8 */
            {8'h00}, /* 0xedb7 */
            {8'h00}, /* 0xedb6 */
            {8'h00}, /* 0xedb5 */
            {8'h00}, /* 0xedb4 */
            {8'h00}, /* 0xedb3 */
            {8'h00}, /* 0xedb2 */
            {8'h00}, /* 0xedb1 */
            {8'h00}, /* 0xedb0 */
            {8'h00}, /* 0xedaf */
            {8'h00}, /* 0xedae */
            {8'h00}, /* 0xedad */
            {8'h00}, /* 0xedac */
            {8'h00}, /* 0xedab */
            {8'h00}, /* 0xedaa */
            {8'h00}, /* 0xeda9 */
            {8'h00}, /* 0xeda8 */
            {8'h00}, /* 0xeda7 */
            {8'h00}, /* 0xeda6 */
            {8'h00}, /* 0xeda5 */
            {8'h00}, /* 0xeda4 */
            {8'h00}, /* 0xeda3 */
            {8'h00}, /* 0xeda2 */
            {8'h00}, /* 0xeda1 */
            {8'h00}, /* 0xeda0 */
            {8'h00}, /* 0xed9f */
            {8'h00}, /* 0xed9e */
            {8'h00}, /* 0xed9d */
            {8'h00}, /* 0xed9c */
            {8'h00}, /* 0xed9b */
            {8'h00}, /* 0xed9a */
            {8'h00}, /* 0xed99 */
            {8'h00}, /* 0xed98 */
            {8'h00}, /* 0xed97 */
            {8'h00}, /* 0xed96 */
            {8'h00}, /* 0xed95 */
            {8'h00}, /* 0xed94 */
            {8'h00}, /* 0xed93 */
            {8'h00}, /* 0xed92 */
            {8'h00}, /* 0xed91 */
            {8'h00}, /* 0xed90 */
            {8'h00}, /* 0xed8f */
            {8'h00}, /* 0xed8e */
            {8'h00}, /* 0xed8d */
            {8'h00}, /* 0xed8c */
            {8'h00}, /* 0xed8b */
            {8'h00}, /* 0xed8a */
            {8'h00}, /* 0xed89 */
            {8'h00}, /* 0xed88 */
            {8'h00}, /* 0xed87 */
            {8'h00}, /* 0xed86 */
            {8'h00}, /* 0xed85 */
            {8'h00}, /* 0xed84 */
            {8'h00}, /* 0xed83 */
            {8'h00}, /* 0xed82 */
            {8'h00}, /* 0xed81 */
            {8'h00}, /* 0xed80 */
            {8'h00}, /* 0xed7f */
            {8'h00}, /* 0xed7e */
            {8'h00}, /* 0xed7d */
            {8'h00}, /* 0xed7c */
            {8'h00}, /* 0xed7b */
            {8'h00}, /* 0xed7a */
            {8'h00}, /* 0xed79 */
            {8'h00}, /* 0xed78 */
            {8'h00}, /* 0xed77 */
            {8'h00}, /* 0xed76 */
            {8'h00}, /* 0xed75 */
            {8'h00}, /* 0xed74 */
            {8'h00}, /* 0xed73 */
            {8'h00}, /* 0xed72 */
            {8'h00}, /* 0xed71 */
            {8'h00}, /* 0xed70 */
            {8'h00}, /* 0xed6f */
            {8'h00}, /* 0xed6e */
            {8'h00}, /* 0xed6d */
            {8'h00}, /* 0xed6c */
            {8'h00}, /* 0xed6b */
            {8'h00}, /* 0xed6a */
            {8'h00}, /* 0xed69 */
            {8'h00}, /* 0xed68 */
            {8'h00}, /* 0xed67 */
            {8'h00}, /* 0xed66 */
            {8'h00}, /* 0xed65 */
            {8'h00}, /* 0xed64 */
            {8'h00}, /* 0xed63 */
            {8'h00}, /* 0xed62 */
            {8'h00}, /* 0xed61 */
            {8'h00}, /* 0xed60 */
            {8'h00}, /* 0xed5f */
            {8'h00}, /* 0xed5e */
            {8'h00}, /* 0xed5d */
            {8'h00}, /* 0xed5c */
            {8'h00}, /* 0xed5b */
            {8'h00}, /* 0xed5a */
            {8'h00}, /* 0xed59 */
            {8'h00}, /* 0xed58 */
            {8'h00}, /* 0xed57 */
            {8'h00}, /* 0xed56 */
            {8'h00}, /* 0xed55 */
            {8'h00}, /* 0xed54 */
            {8'h00}, /* 0xed53 */
            {8'h00}, /* 0xed52 */
            {8'h00}, /* 0xed51 */
            {8'h00}, /* 0xed50 */
            {8'h00}, /* 0xed4f */
            {8'h00}, /* 0xed4e */
            {8'h00}, /* 0xed4d */
            {8'h00}, /* 0xed4c */
            {8'h00}, /* 0xed4b */
            {8'h00}, /* 0xed4a */
            {8'h00}, /* 0xed49 */
            {8'h00}, /* 0xed48 */
            {8'h00}, /* 0xed47 */
            {8'h00}, /* 0xed46 */
            {8'h00}, /* 0xed45 */
            {8'h00}, /* 0xed44 */
            {8'h00}, /* 0xed43 */
            {8'h00}, /* 0xed42 */
            {8'h00}, /* 0xed41 */
            {8'h00}, /* 0xed40 */
            {8'h00}, /* 0xed3f */
            {8'h00}, /* 0xed3e */
            {8'h00}, /* 0xed3d */
            {8'h00}, /* 0xed3c */
            {8'h00}, /* 0xed3b */
            {8'h00}, /* 0xed3a */
            {8'h00}, /* 0xed39 */
            {8'h00}, /* 0xed38 */
            {8'h00}, /* 0xed37 */
            {8'h00}, /* 0xed36 */
            {8'h00}, /* 0xed35 */
            {8'h00}, /* 0xed34 */
            {8'h00}, /* 0xed33 */
            {8'h00}, /* 0xed32 */
            {8'h00}, /* 0xed31 */
            {8'h00}, /* 0xed30 */
            {8'h00}, /* 0xed2f */
            {8'h00}, /* 0xed2e */
            {8'h00}, /* 0xed2d */
            {8'h00}, /* 0xed2c */
            {8'h00}, /* 0xed2b */
            {8'h00}, /* 0xed2a */
            {8'h00}, /* 0xed29 */
            {8'h00}, /* 0xed28 */
            {8'h00}, /* 0xed27 */
            {8'h00}, /* 0xed26 */
            {8'h00}, /* 0xed25 */
            {8'h00}, /* 0xed24 */
            {8'h00}, /* 0xed23 */
            {8'h00}, /* 0xed22 */
            {8'h00}, /* 0xed21 */
            {8'h00}, /* 0xed20 */
            {8'h00}, /* 0xed1f */
            {8'h00}, /* 0xed1e */
            {8'h00}, /* 0xed1d */
            {8'h00}, /* 0xed1c */
            {8'h00}, /* 0xed1b */
            {8'h00}, /* 0xed1a */
            {8'h00}, /* 0xed19 */
            {8'h00}, /* 0xed18 */
            {8'h00}, /* 0xed17 */
            {8'h00}, /* 0xed16 */
            {8'h00}, /* 0xed15 */
            {8'h00}, /* 0xed14 */
            {8'h00}, /* 0xed13 */
            {8'h00}, /* 0xed12 */
            {8'h00}, /* 0xed11 */
            {8'h00}, /* 0xed10 */
            {8'h00}, /* 0xed0f */
            {8'h00}, /* 0xed0e */
            {8'h00}, /* 0xed0d */
            {8'h00}, /* 0xed0c */
            {8'h00}, /* 0xed0b */
            {8'h00}, /* 0xed0a */
            {8'h00}, /* 0xed09 */
            {8'h00}, /* 0xed08 */
            {8'h00}, /* 0xed07 */
            {8'h00}, /* 0xed06 */
            {8'h00}, /* 0xed05 */
            {8'h00}, /* 0xed04 */
            {8'h00}, /* 0xed03 */
            {8'h00}, /* 0xed02 */
            {8'h00}, /* 0xed01 */
            {8'h00}, /* 0xed00 */
            {8'h00}, /* 0xecff */
            {8'h00}, /* 0xecfe */
            {8'h00}, /* 0xecfd */
            {8'h00}, /* 0xecfc */
            {8'h00}, /* 0xecfb */
            {8'h00}, /* 0xecfa */
            {8'h00}, /* 0xecf9 */
            {8'h00}, /* 0xecf8 */
            {8'h00}, /* 0xecf7 */
            {8'h00}, /* 0xecf6 */
            {8'h00}, /* 0xecf5 */
            {8'h00}, /* 0xecf4 */
            {8'h00}, /* 0xecf3 */
            {8'h00}, /* 0xecf2 */
            {8'h00}, /* 0xecf1 */
            {8'h00}, /* 0xecf0 */
            {8'h00}, /* 0xecef */
            {8'h00}, /* 0xecee */
            {8'h00}, /* 0xeced */
            {8'h00}, /* 0xecec */
            {8'h00}, /* 0xeceb */
            {8'h00}, /* 0xecea */
            {8'h00}, /* 0xece9 */
            {8'h00}, /* 0xece8 */
            {8'h00}, /* 0xece7 */
            {8'h00}, /* 0xece6 */
            {8'h00}, /* 0xece5 */
            {8'h00}, /* 0xece4 */
            {8'h00}, /* 0xece3 */
            {8'h00}, /* 0xece2 */
            {8'h00}, /* 0xece1 */
            {8'h00}, /* 0xece0 */
            {8'h00}, /* 0xecdf */
            {8'h00}, /* 0xecde */
            {8'h00}, /* 0xecdd */
            {8'h00}, /* 0xecdc */
            {8'h00}, /* 0xecdb */
            {8'h00}, /* 0xecda */
            {8'h00}, /* 0xecd9 */
            {8'h00}, /* 0xecd8 */
            {8'h00}, /* 0xecd7 */
            {8'h00}, /* 0xecd6 */
            {8'h00}, /* 0xecd5 */
            {8'h00}, /* 0xecd4 */
            {8'h00}, /* 0xecd3 */
            {8'h00}, /* 0xecd2 */
            {8'h00}, /* 0xecd1 */
            {8'h00}, /* 0xecd0 */
            {8'h00}, /* 0xeccf */
            {8'h00}, /* 0xecce */
            {8'h00}, /* 0xeccd */
            {8'h00}, /* 0xeccc */
            {8'h00}, /* 0xeccb */
            {8'h00}, /* 0xecca */
            {8'h00}, /* 0xecc9 */
            {8'h00}, /* 0xecc8 */
            {8'h00}, /* 0xecc7 */
            {8'h00}, /* 0xecc6 */
            {8'h00}, /* 0xecc5 */
            {8'h00}, /* 0xecc4 */
            {8'h00}, /* 0xecc3 */
            {8'h00}, /* 0xecc2 */
            {8'h00}, /* 0xecc1 */
            {8'h00}, /* 0xecc0 */
            {8'h00}, /* 0xecbf */
            {8'h00}, /* 0xecbe */
            {8'h00}, /* 0xecbd */
            {8'h00}, /* 0xecbc */
            {8'h00}, /* 0xecbb */
            {8'h00}, /* 0xecba */
            {8'h00}, /* 0xecb9 */
            {8'h00}, /* 0xecb8 */
            {8'h00}, /* 0xecb7 */
            {8'h00}, /* 0xecb6 */
            {8'h00}, /* 0xecb5 */
            {8'h00}, /* 0xecb4 */
            {8'h00}, /* 0xecb3 */
            {8'h00}, /* 0xecb2 */
            {8'h00}, /* 0xecb1 */
            {8'h00}, /* 0xecb0 */
            {8'h00}, /* 0xecaf */
            {8'h00}, /* 0xecae */
            {8'h00}, /* 0xecad */
            {8'h00}, /* 0xecac */
            {8'h00}, /* 0xecab */
            {8'h00}, /* 0xecaa */
            {8'h00}, /* 0xeca9 */
            {8'h00}, /* 0xeca8 */
            {8'h00}, /* 0xeca7 */
            {8'h00}, /* 0xeca6 */
            {8'h00}, /* 0xeca5 */
            {8'h00}, /* 0xeca4 */
            {8'h00}, /* 0xeca3 */
            {8'h00}, /* 0xeca2 */
            {8'h00}, /* 0xeca1 */
            {8'h00}, /* 0xeca0 */
            {8'h00}, /* 0xec9f */
            {8'h00}, /* 0xec9e */
            {8'h00}, /* 0xec9d */
            {8'h00}, /* 0xec9c */
            {8'h00}, /* 0xec9b */
            {8'h00}, /* 0xec9a */
            {8'h00}, /* 0xec99 */
            {8'h00}, /* 0xec98 */
            {8'h00}, /* 0xec97 */
            {8'h00}, /* 0xec96 */
            {8'h00}, /* 0xec95 */
            {8'h00}, /* 0xec94 */
            {8'h00}, /* 0xec93 */
            {8'h00}, /* 0xec92 */
            {8'h00}, /* 0xec91 */
            {8'h00}, /* 0xec90 */
            {8'h00}, /* 0xec8f */
            {8'h00}, /* 0xec8e */
            {8'h00}, /* 0xec8d */
            {8'h00}, /* 0xec8c */
            {8'h00}, /* 0xec8b */
            {8'h00}, /* 0xec8a */
            {8'h00}, /* 0xec89 */
            {8'h00}, /* 0xec88 */
            {8'h00}, /* 0xec87 */
            {8'h00}, /* 0xec86 */
            {8'h00}, /* 0xec85 */
            {8'h00}, /* 0xec84 */
            {8'h00}, /* 0xec83 */
            {8'h00}, /* 0xec82 */
            {8'h00}, /* 0xec81 */
            {8'h00}, /* 0xec80 */
            {8'h00}, /* 0xec7f */
            {8'h00}, /* 0xec7e */
            {8'h00}, /* 0xec7d */
            {8'h00}, /* 0xec7c */
            {8'h00}, /* 0xec7b */
            {8'h00}, /* 0xec7a */
            {8'h00}, /* 0xec79 */
            {8'h00}, /* 0xec78 */
            {8'h00}, /* 0xec77 */
            {8'h00}, /* 0xec76 */
            {8'h00}, /* 0xec75 */
            {8'h00}, /* 0xec74 */
            {8'h00}, /* 0xec73 */
            {8'h00}, /* 0xec72 */
            {8'h00}, /* 0xec71 */
            {8'h00}, /* 0xec70 */
            {8'h00}, /* 0xec6f */
            {8'h00}, /* 0xec6e */
            {8'h00}, /* 0xec6d */
            {8'h00}, /* 0xec6c */
            {8'h00}, /* 0xec6b */
            {8'h00}, /* 0xec6a */
            {8'h00}, /* 0xec69 */
            {8'h00}, /* 0xec68 */
            {8'h00}, /* 0xec67 */
            {8'h00}, /* 0xec66 */
            {8'h00}, /* 0xec65 */
            {8'h00}, /* 0xec64 */
            {8'h00}, /* 0xec63 */
            {8'h00}, /* 0xec62 */
            {8'h00}, /* 0xec61 */
            {8'h00}, /* 0xec60 */
            {8'h00}, /* 0xec5f */
            {8'h00}, /* 0xec5e */
            {8'h00}, /* 0xec5d */
            {8'h00}, /* 0xec5c */
            {8'h00}, /* 0xec5b */
            {8'h00}, /* 0xec5a */
            {8'h00}, /* 0xec59 */
            {8'h00}, /* 0xec58 */
            {8'h00}, /* 0xec57 */
            {8'h00}, /* 0xec56 */
            {8'h00}, /* 0xec55 */
            {8'h00}, /* 0xec54 */
            {8'h00}, /* 0xec53 */
            {8'h00}, /* 0xec52 */
            {8'h00}, /* 0xec51 */
            {8'h00}, /* 0xec50 */
            {8'h00}, /* 0xec4f */
            {8'h00}, /* 0xec4e */
            {8'h00}, /* 0xec4d */
            {8'h00}, /* 0xec4c */
            {8'h00}, /* 0xec4b */
            {8'h00}, /* 0xec4a */
            {8'h00}, /* 0xec49 */
            {8'h00}, /* 0xec48 */
            {8'h00}, /* 0xec47 */
            {8'h00}, /* 0xec46 */
            {8'h00}, /* 0xec45 */
            {8'h00}, /* 0xec44 */
            {8'h00}, /* 0xec43 */
            {8'h00}, /* 0xec42 */
            {8'h00}, /* 0xec41 */
            {8'h00}, /* 0xec40 */
            {8'h00}, /* 0xec3f */
            {8'h00}, /* 0xec3e */
            {8'h00}, /* 0xec3d */
            {8'h00}, /* 0xec3c */
            {8'h00}, /* 0xec3b */
            {8'h00}, /* 0xec3a */
            {8'h00}, /* 0xec39 */
            {8'h00}, /* 0xec38 */
            {8'h00}, /* 0xec37 */
            {8'h00}, /* 0xec36 */
            {8'h00}, /* 0xec35 */
            {8'h00}, /* 0xec34 */
            {8'h00}, /* 0xec33 */
            {8'h00}, /* 0xec32 */
            {8'h00}, /* 0xec31 */
            {8'h00}, /* 0xec30 */
            {8'h00}, /* 0xec2f */
            {8'h00}, /* 0xec2e */
            {8'h00}, /* 0xec2d */
            {8'h00}, /* 0xec2c */
            {8'h00}, /* 0xec2b */
            {8'h00}, /* 0xec2a */
            {8'h00}, /* 0xec29 */
            {8'h00}, /* 0xec28 */
            {8'h00}, /* 0xec27 */
            {8'h00}, /* 0xec26 */
            {8'h00}, /* 0xec25 */
            {8'h00}, /* 0xec24 */
            {8'h00}, /* 0xec23 */
            {8'h00}, /* 0xec22 */
            {8'h00}, /* 0xec21 */
            {8'h00}, /* 0xec20 */
            {8'h00}, /* 0xec1f */
            {8'h00}, /* 0xec1e */
            {8'h00}, /* 0xec1d */
            {8'h00}, /* 0xec1c */
            {8'h00}, /* 0xec1b */
            {8'h00}, /* 0xec1a */
            {8'h00}, /* 0xec19 */
            {8'h00}, /* 0xec18 */
            {8'h00}, /* 0xec17 */
            {8'h00}, /* 0xec16 */
            {8'h00}, /* 0xec15 */
            {8'h00}, /* 0xec14 */
            {8'h00}, /* 0xec13 */
            {8'h00}, /* 0xec12 */
            {8'h00}, /* 0xec11 */
            {8'h00}, /* 0xec10 */
            {8'h00}, /* 0xec0f */
            {8'h00}, /* 0xec0e */
            {8'h00}, /* 0xec0d */
            {8'h00}, /* 0xec0c */
            {8'h00}, /* 0xec0b */
            {8'h00}, /* 0xec0a */
            {8'h00}, /* 0xec09 */
            {8'h00}, /* 0xec08 */
            {8'h00}, /* 0xec07 */
            {8'h00}, /* 0xec06 */
            {8'h00}, /* 0xec05 */
            {8'h00}, /* 0xec04 */
            {8'h00}, /* 0xec03 */
            {8'h00}, /* 0xec02 */
            {8'h00}, /* 0xec01 */
            {8'h00}, /* 0xec00 */
            {8'h00}, /* 0xebff */
            {8'h00}, /* 0xebfe */
            {8'h00}, /* 0xebfd */
            {8'h00}, /* 0xebfc */
            {8'h00}, /* 0xebfb */
            {8'h00}, /* 0xebfa */
            {8'h00}, /* 0xebf9 */
            {8'h00}, /* 0xebf8 */
            {8'h00}, /* 0xebf7 */
            {8'h00}, /* 0xebf6 */
            {8'h00}, /* 0xebf5 */
            {8'h00}, /* 0xebf4 */
            {8'h00}, /* 0xebf3 */
            {8'h00}, /* 0xebf2 */
            {8'h00}, /* 0xebf1 */
            {8'h00}, /* 0xebf0 */
            {8'h00}, /* 0xebef */
            {8'h00}, /* 0xebee */
            {8'h00}, /* 0xebed */
            {8'h00}, /* 0xebec */
            {8'h00}, /* 0xebeb */
            {8'h00}, /* 0xebea */
            {8'h00}, /* 0xebe9 */
            {8'h00}, /* 0xebe8 */
            {8'h00}, /* 0xebe7 */
            {8'h00}, /* 0xebe6 */
            {8'h00}, /* 0xebe5 */
            {8'h00}, /* 0xebe4 */
            {8'h00}, /* 0xebe3 */
            {8'h00}, /* 0xebe2 */
            {8'h00}, /* 0xebe1 */
            {8'h00}, /* 0xebe0 */
            {8'h00}, /* 0xebdf */
            {8'h00}, /* 0xebde */
            {8'h00}, /* 0xebdd */
            {8'h00}, /* 0xebdc */
            {8'h00}, /* 0xebdb */
            {8'h00}, /* 0xebda */
            {8'h00}, /* 0xebd9 */
            {8'h00}, /* 0xebd8 */
            {8'h00}, /* 0xebd7 */
            {8'h00}, /* 0xebd6 */
            {8'h00}, /* 0xebd5 */
            {8'h00}, /* 0xebd4 */
            {8'h00}, /* 0xebd3 */
            {8'h00}, /* 0xebd2 */
            {8'h00}, /* 0xebd1 */
            {8'h00}, /* 0xebd0 */
            {8'h00}, /* 0xebcf */
            {8'h00}, /* 0xebce */
            {8'h00}, /* 0xebcd */
            {8'h00}, /* 0xebcc */
            {8'h00}, /* 0xebcb */
            {8'h00}, /* 0xebca */
            {8'h00}, /* 0xebc9 */
            {8'h00}, /* 0xebc8 */
            {8'h00}, /* 0xebc7 */
            {8'h00}, /* 0xebc6 */
            {8'h00}, /* 0xebc5 */
            {8'h00}, /* 0xebc4 */
            {8'h00}, /* 0xebc3 */
            {8'h00}, /* 0xebc2 */
            {8'h00}, /* 0xebc1 */
            {8'h00}, /* 0xebc0 */
            {8'h00}, /* 0xebbf */
            {8'h00}, /* 0xebbe */
            {8'h00}, /* 0xebbd */
            {8'h00}, /* 0xebbc */
            {8'h00}, /* 0xebbb */
            {8'h00}, /* 0xebba */
            {8'h00}, /* 0xebb9 */
            {8'h00}, /* 0xebb8 */
            {8'h00}, /* 0xebb7 */
            {8'h00}, /* 0xebb6 */
            {8'h00}, /* 0xebb5 */
            {8'h00}, /* 0xebb4 */
            {8'h00}, /* 0xebb3 */
            {8'h00}, /* 0xebb2 */
            {8'h00}, /* 0xebb1 */
            {8'h00}, /* 0xebb0 */
            {8'h00}, /* 0xebaf */
            {8'h00}, /* 0xebae */
            {8'h00}, /* 0xebad */
            {8'h00}, /* 0xebac */
            {8'h00}, /* 0xebab */
            {8'h00}, /* 0xebaa */
            {8'h00}, /* 0xeba9 */
            {8'h00}, /* 0xeba8 */
            {8'h00}, /* 0xeba7 */
            {8'h00}, /* 0xeba6 */
            {8'h00}, /* 0xeba5 */
            {8'h00}, /* 0xeba4 */
            {8'h00}, /* 0xeba3 */
            {8'h00}, /* 0xeba2 */
            {8'h00}, /* 0xeba1 */
            {8'h00}, /* 0xeba0 */
            {8'h00}, /* 0xeb9f */
            {8'h00}, /* 0xeb9e */
            {8'h00}, /* 0xeb9d */
            {8'h00}, /* 0xeb9c */
            {8'h00}, /* 0xeb9b */
            {8'h00}, /* 0xeb9a */
            {8'h00}, /* 0xeb99 */
            {8'h00}, /* 0xeb98 */
            {8'h00}, /* 0xeb97 */
            {8'h00}, /* 0xeb96 */
            {8'h00}, /* 0xeb95 */
            {8'h00}, /* 0xeb94 */
            {8'h00}, /* 0xeb93 */
            {8'h00}, /* 0xeb92 */
            {8'h00}, /* 0xeb91 */
            {8'h00}, /* 0xeb90 */
            {8'h00}, /* 0xeb8f */
            {8'h00}, /* 0xeb8e */
            {8'h00}, /* 0xeb8d */
            {8'h00}, /* 0xeb8c */
            {8'h00}, /* 0xeb8b */
            {8'h00}, /* 0xeb8a */
            {8'h00}, /* 0xeb89 */
            {8'h00}, /* 0xeb88 */
            {8'h00}, /* 0xeb87 */
            {8'h00}, /* 0xeb86 */
            {8'h00}, /* 0xeb85 */
            {8'h00}, /* 0xeb84 */
            {8'h00}, /* 0xeb83 */
            {8'h00}, /* 0xeb82 */
            {8'h00}, /* 0xeb81 */
            {8'h00}, /* 0xeb80 */
            {8'h00}, /* 0xeb7f */
            {8'h00}, /* 0xeb7e */
            {8'h00}, /* 0xeb7d */
            {8'h00}, /* 0xeb7c */
            {8'h00}, /* 0xeb7b */
            {8'h00}, /* 0xeb7a */
            {8'h00}, /* 0xeb79 */
            {8'h00}, /* 0xeb78 */
            {8'h00}, /* 0xeb77 */
            {8'h00}, /* 0xeb76 */
            {8'h00}, /* 0xeb75 */
            {8'h00}, /* 0xeb74 */
            {8'h00}, /* 0xeb73 */
            {8'h00}, /* 0xeb72 */
            {8'h00}, /* 0xeb71 */
            {8'h00}, /* 0xeb70 */
            {8'h00}, /* 0xeb6f */
            {8'h00}, /* 0xeb6e */
            {8'h00}, /* 0xeb6d */
            {8'h00}, /* 0xeb6c */
            {8'h00}, /* 0xeb6b */
            {8'h00}, /* 0xeb6a */
            {8'h00}, /* 0xeb69 */
            {8'h00}, /* 0xeb68 */
            {8'h00}, /* 0xeb67 */
            {8'h00}, /* 0xeb66 */
            {8'h00}, /* 0xeb65 */
            {8'h00}, /* 0xeb64 */
            {8'h00}, /* 0xeb63 */
            {8'h00}, /* 0xeb62 */
            {8'h00}, /* 0xeb61 */
            {8'h00}, /* 0xeb60 */
            {8'h00}, /* 0xeb5f */
            {8'h00}, /* 0xeb5e */
            {8'h00}, /* 0xeb5d */
            {8'h00}, /* 0xeb5c */
            {8'h00}, /* 0xeb5b */
            {8'h00}, /* 0xeb5a */
            {8'h00}, /* 0xeb59 */
            {8'h00}, /* 0xeb58 */
            {8'h00}, /* 0xeb57 */
            {8'h00}, /* 0xeb56 */
            {8'h00}, /* 0xeb55 */
            {8'h00}, /* 0xeb54 */
            {8'h00}, /* 0xeb53 */
            {8'h00}, /* 0xeb52 */
            {8'h00}, /* 0xeb51 */
            {8'h00}, /* 0xeb50 */
            {8'h00}, /* 0xeb4f */
            {8'h00}, /* 0xeb4e */
            {8'h00}, /* 0xeb4d */
            {8'h00}, /* 0xeb4c */
            {8'h00}, /* 0xeb4b */
            {8'h00}, /* 0xeb4a */
            {8'h00}, /* 0xeb49 */
            {8'h00}, /* 0xeb48 */
            {8'h00}, /* 0xeb47 */
            {8'h00}, /* 0xeb46 */
            {8'h00}, /* 0xeb45 */
            {8'h00}, /* 0xeb44 */
            {8'h00}, /* 0xeb43 */
            {8'h00}, /* 0xeb42 */
            {8'h00}, /* 0xeb41 */
            {8'h00}, /* 0xeb40 */
            {8'h00}, /* 0xeb3f */
            {8'h00}, /* 0xeb3e */
            {8'h00}, /* 0xeb3d */
            {8'h00}, /* 0xeb3c */
            {8'h00}, /* 0xeb3b */
            {8'h00}, /* 0xeb3a */
            {8'h00}, /* 0xeb39 */
            {8'h00}, /* 0xeb38 */
            {8'h00}, /* 0xeb37 */
            {8'h00}, /* 0xeb36 */
            {8'h00}, /* 0xeb35 */
            {8'h00}, /* 0xeb34 */
            {8'h00}, /* 0xeb33 */
            {8'h00}, /* 0xeb32 */
            {8'h00}, /* 0xeb31 */
            {8'h00}, /* 0xeb30 */
            {8'h00}, /* 0xeb2f */
            {8'h00}, /* 0xeb2e */
            {8'h00}, /* 0xeb2d */
            {8'h00}, /* 0xeb2c */
            {8'h00}, /* 0xeb2b */
            {8'h00}, /* 0xeb2a */
            {8'h00}, /* 0xeb29 */
            {8'h00}, /* 0xeb28 */
            {8'h00}, /* 0xeb27 */
            {8'h00}, /* 0xeb26 */
            {8'h00}, /* 0xeb25 */
            {8'h00}, /* 0xeb24 */
            {8'h00}, /* 0xeb23 */
            {8'h00}, /* 0xeb22 */
            {8'h00}, /* 0xeb21 */
            {8'h00}, /* 0xeb20 */
            {8'h00}, /* 0xeb1f */
            {8'h00}, /* 0xeb1e */
            {8'h00}, /* 0xeb1d */
            {8'h00}, /* 0xeb1c */
            {8'h00}, /* 0xeb1b */
            {8'h00}, /* 0xeb1a */
            {8'h00}, /* 0xeb19 */
            {8'h00}, /* 0xeb18 */
            {8'h00}, /* 0xeb17 */
            {8'h00}, /* 0xeb16 */
            {8'h00}, /* 0xeb15 */
            {8'h00}, /* 0xeb14 */
            {8'h00}, /* 0xeb13 */
            {8'h00}, /* 0xeb12 */
            {8'h00}, /* 0xeb11 */
            {8'h00}, /* 0xeb10 */
            {8'h00}, /* 0xeb0f */
            {8'h00}, /* 0xeb0e */
            {8'h00}, /* 0xeb0d */
            {8'h00}, /* 0xeb0c */
            {8'h00}, /* 0xeb0b */
            {8'h00}, /* 0xeb0a */
            {8'h00}, /* 0xeb09 */
            {8'h00}, /* 0xeb08 */
            {8'h00}, /* 0xeb07 */
            {8'h00}, /* 0xeb06 */
            {8'h00}, /* 0xeb05 */
            {8'h00}, /* 0xeb04 */
            {8'h00}, /* 0xeb03 */
            {8'h00}, /* 0xeb02 */
            {8'h00}, /* 0xeb01 */
            {8'h00}, /* 0xeb00 */
            {8'h00}, /* 0xeaff */
            {8'h00}, /* 0xeafe */
            {8'h00}, /* 0xeafd */
            {8'h00}, /* 0xeafc */
            {8'h00}, /* 0xeafb */
            {8'h00}, /* 0xeafa */
            {8'h00}, /* 0xeaf9 */
            {8'h00}, /* 0xeaf8 */
            {8'h00}, /* 0xeaf7 */
            {8'h00}, /* 0xeaf6 */
            {8'h00}, /* 0xeaf5 */
            {8'h00}, /* 0xeaf4 */
            {8'h00}, /* 0xeaf3 */
            {8'h00}, /* 0xeaf2 */
            {8'h00}, /* 0xeaf1 */
            {8'h00}, /* 0xeaf0 */
            {8'h00}, /* 0xeaef */
            {8'h00}, /* 0xeaee */
            {8'h00}, /* 0xeaed */
            {8'h00}, /* 0xeaec */
            {8'h00}, /* 0xeaeb */
            {8'h00}, /* 0xeaea */
            {8'h00}, /* 0xeae9 */
            {8'h00}, /* 0xeae8 */
            {8'h00}, /* 0xeae7 */
            {8'h00}, /* 0xeae6 */
            {8'h00}, /* 0xeae5 */
            {8'h00}, /* 0xeae4 */
            {8'h00}, /* 0xeae3 */
            {8'h00}, /* 0xeae2 */
            {8'h00}, /* 0xeae1 */
            {8'h00}, /* 0xeae0 */
            {8'h00}, /* 0xeadf */
            {8'h00}, /* 0xeade */
            {8'h00}, /* 0xeadd */
            {8'h00}, /* 0xeadc */
            {8'h00}, /* 0xeadb */
            {8'h00}, /* 0xeada */
            {8'h00}, /* 0xead9 */
            {8'h00}, /* 0xead8 */
            {8'h00}, /* 0xead7 */
            {8'h00}, /* 0xead6 */
            {8'h00}, /* 0xead5 */
            {8'h00}, /* 0xead4 */
            {8'h00}, /* 0xead3 */
            {8'h00}, /* 0xead2 */
            {8'h00}, /* 0xead1 */
            {8'h00}, /* 0xead0 */
            {8'h00}, /* 0xeacf */
            {8'h00}, /* 0xeace */
            {8'h00}, /* 0xeacd */
            {8'h00}, /* 0xeacc */
            {8'h00}, /* 0xeacb */
            {8'h00}, /* 0xeaca */
            {8'h00}, /* 0xeac9 */
            {8'h00}, /* 0xeac8 */
            {8'h00}, /* 0xeac7 */
            {8'h00}, /* 0xeac6 */
            {8'h00}, /* 0xeac5 */
            {8'h00}, /* 0xeac4 */
            {8'h00}, /* 0xeac3 */
            {8'h00}, /* 0xeac2 */
            {8'h00}, /* 0xeac1 */
            {8'h00}, /* 0xeac0 */
            {8'h00}, /* 0xeabf */
            {8'h00}, /* 0xeabe */
            {8'h00}, /* 0xeabd */
            {8'h00}, /* 0xeabc */
            {8'h00}, /* 0xeabb */
            {8'h00}, /* 0xeaba */
            {8'h00}, /* 0xeab9 */
            {8'h00}, /* 0xeab8 */
            {8'h00}, /* 0xeab7 */
            {8'h00}, /* 0xeab6 */
            {8'h00}, /* 0xeab5 */
            {8'h00}, /* 0xeab4 */
            {8'h00}, /* 0xeab3 */
            {8'h00}, /* 0xeab2 */
            {8'h00}, /* 0xeab1 */
            {8'h00}, /* 0xeab0 */
            {8'h00}, /* 0xeaaf */
            {8'h00}, /* 0xeaae */
            {8'h00}, /* 0xeaad */
            {8'h00}, /* 0xeaac */
            {8'h00}, /* 0xeaab */
            {8'h00}, /* 0xeaaa */
            {8'h00}, /* 0xeaa9 */
            {8'h00}, /* 0xeaa8 */
            {8'h00}, /* 0xeaa7 */
            {8'h00}, /* 0xeaa6 */
            {8'h00}, /* 0xeaa5 */
            {8'h00}, /* 0xeaa4 */
            {8'h00}, /* 0xeaa3 */
            {8'h00}, /* 0xeaa2 */
            {8'h00}, /* 0xeaa1 */
            {8'h00}, /* 0xeaa0 */
            {8'h00}, /* 0xea9f */
            {8'h00}, /* 0xea9e */
            {8'h00}, /* 0xea9d */
            {8'h00}, /* 0xea9c */
            {8'h00}, /* 0xea9b */
            {8'h00}, /* 0xea9a */
            {8'h00}, /* 0xea99 */
            {8'h00}, /* 0xea98 */
            {8'h00}, /* 0xea97 */
            {8'h00}, /* 0xea96 */
            {8'h00}, /* 0xea95 */
            {8'h00}, /* 0xea94 */
            {8'h00}, /* 0xea93 */
            {8'h00}, /* 0xea92 */
            {8'h00}, /* 0xea91 */
            {8'h00}, /* 0xea90 */
            {8'h00}, /* 0xea8f */
            {8'h00}, /* 0xea8e */
            {8'h00}, /* 0xea8d */
            {8'h00}, /* 0xea8c */
            {8'h00}, /* 0xea8b */
            {8'h00}, /* 0xea8a */
            {8'h00}, /* 0xea89 */
            {8'h00}, /* 0xea88 */
            {8'h00}, /* 0xea87 */
            {8'h00}, /* 0xea86 */
            {8'h00}, /* 0xea85 */
            {8'h00}, /* 0xea84 */
            {8'h00}, /* 0xea83 */
            {8'h00}, /* 0xea82 */
            {8'h00}, /* 0xea81 */
            {8'h00}, /* 0xea80 */
            {8'h00}, /* 0xea7f */
            {8'h00}, /* 0xea7e */
            {8'h00}, /* 0xea7d */
            {8'h00}, /* 0xea7c */
            {8'h00}, /* 0xea7b */
            {8'h00}, /* 0xea7a */
            {8'h00}, /* 0xea79 */
            {8'h00}, /* 0xea78 */
            {8'h00}, /* 0xea77 */
            {8'h00}, /* 0xea76 */
            {8'h00}, /* 0xea75 */
            {8'h00}, /* 0xea74 */
            {8'h00}, /* 0xea73 */
            {8'h00}, /* 0xea72 */
            {8'h00}, /* 0xea71 */
            {8'h00}, /* 0xea70 */
            {8'h00}, /* 0xea6f */
            {8'h00}, /* 0xea6e */
            {8'h00}, /* 0xea6d */
            {8'h00}, /* 0xea6c */
            {8'h00}, /* 0xea6b */
            {8'h00}, /* 0xea6a */
            {8'h00}, /* 0xea69 */
            {8'h00}, /* 0xea68 */
            {8'h00}, /* 0xea67 */
            {8'h00}, /* 0xea66 */
            {8'h00}, /* 0xea65 */
            {8'h00}, /* 0xea64 */
            {8'h00}, /* 0xea63 */
            {8'h00}, /* 0xea62 */
            {8'h00}, /* 0xea61 */
            {8'h00}, /* 0xea60 */
            {8'h00}, /* 0xea5f */
            {8'h00}, /* 0xea5e */
            {8'h00}, /* 0xea5d */
            {8'h00}, /* 0xea5c */
            {8'h00}, /* 0xea5b */
            {8'h00}, /* 0xea5a */
            {8'h00}, /* 0xea59 */
            {8'h00}, /* 0xea58 */
            {8'h00}, /* 0xea57 */
            {8'h00}, /* 0xea56 */
            {8'h00}, /* 0xea55 */
            {8'h00}, /* 0xea54 */
            {8'h00}, /* 0xea53 */
            {8'h00}, /* 0xea52 */
            {8'h00}, /* 0xea51 */
            {8'h00}, /* 0xea50 */
            {8'h00}, /* 0xea4f */
            {8'h00}, /* 0xea4e */
            {8'h00}, /* 0xea4d */
            {8'h00}, /* 0xea4c */
            {8'h00}, /* 0xea4b */
            {8'h00}, /* 0xea4a */
            {8'h00}, /* 0xea49 */
            {8'h00}, /* 0xea48 */
            {8'h00}, /* 0xea47 */
            {8'h00}, /* 0xea46 */
            {8'h00}, /* 0xea45 */
            {8'h00}, /* 0xea44 */
            {8'h00}, /* 0xea43 */
            {8'h00}, /* 0xea42 */
            {8'h00}, /* 0xea41 */
            {8'h00}, /* 0xea40 */
            {8'h00}, /* 0xea3f */
            {8'h00}, /* 0xea3e */
            {8'h00}, /* 0xea3d */
            {8'h00}, /* 0xea3c */
            {8'h00}, /* 0xea3b */
            {8'h00}, /* 0xea3a */
            {8'h00}, /* 0xea39 */
            {8'h00}, /* 0xea38 */
            {8'h00}, /* 0xea37 */
            {8'h00}, /* 0xea36 */
            {8'h00}, /* 0xea35 */
            {8'h00}, /* 0xea34 */
            {8'h00}, /* 0xea33 */
            {8'h00}, /* 0xea32 */
            {8'h00}, /* 0xea31 */
            {8'h00}, /* 0xea30 */
            {8'h00}, /* 0xea2f */
            {8'h00}, /* 0xea2e */
            {8'h00}, /* 0xea2d */
            {8'h00}, /* 0xea2c */
            {8'h00}, /* 0xea2b */
            {8'h00}, /* 0xea2a */
            {8'h00}, /* 0xea29 */
            {8'h00}, /* 0xea28 */
            {8'h00}, /* 0xea27 */
            {8'h00}, /* 0xea26 */
            {8'h00}, /* 0xea25 */
            {8'h00}, /* 0xea24 */
            {8'h00}, /* 0xea23 */
            {8'h00}, /* 0xea22 */
            {8'h00}, /* 0xea21 */
            {8'h00}, /* 0xea20 */
            {8'h00}, /* 0xea1f */
            {8'h00}, /* 0xea1e */
            {8'h00}, /* 0xea1d */
            {8'h00}, /* 0xea1c */
            {8'h00}, /* 0xea1b */
            {8'h00}, /* 0xea1a */
            {8'h00}, /* 0xea19 */
            {8'h00}, /* 0xea18 */
            {8'h00}, /* 0xea17 */
            {8'h00}, /* 0xea16 */
            {8'h00}, /* 0xea15 */
            {8'h00}, /* 0xea14 */
            {8'h00}, /* 0xea13 */
            {8'h00}, /* 0xea12 */
            {8'h00}, /* 0xea11 */
            {8'h00}, /* 0xea10 */
            {8'h00}, /* 0xea0f */
            {8'h00}, /* 0xea0e */
            {8'h00}, /* 0xea0d */
            {8'h00}, /* 0xea0c */
            {8'h00}, /* 0xea0b */
            {8'h00}, /* 0xea0a */
            {8'h00}, /* 0xea09 */
            {8'h00}, /* 0xea08 */
            {8'h00}, /* 0xea07 */
            {8'h00}, /* 0xea06 */
            {8'h00}, /* 0xea05 */
            {8'h00}, /* 0xea04 */
            {8'h00}, /* 0xea03 */
            {8'h00}, /* 0xea02 */
            {8'h00}, /* 0xea01 */
            {8'h00}, /* 0xea00 */
            {8'h00}, /* 0xe9ff */
            {8'h00}, /* 0xe9fe */
            {8'h00}, /* 0xe9fd */
            {8'h00}, /* 0xe9fc */
            {8'h00}, /* 0xe9fb */
            {8'h00}, /* 0xe9fa */
            {8'h00}, /* 0xe9f9 */
            {8'h00}, /* 0xe9f8 */
            {8'h00}, /* 0xe9f7 */
            {8'h00}, /* 0xe9f6 */
            {8'h00}, /* 0xe9f5 */
            {8'h00}, /* 0xe9f4 */
            {8'h00}, /* 0xe9f3 */
            {8'h00}, /* 0xe9f2 */
            {8'h00}, /* 0xe9f1 */
            {8'h00}, /* 0xe9f0 */
            {8'h00}, /* 0xe9ef */
            {8'h00}, /* 0xe9ee */
            {8'h00}, /* 0xe9ed */
            {8'h00}, /* 0xe9ec */
            {8'h00}, /* 0xe9eb */
            {8'h00}, /* 0xe9ea */
            {8'h00}, /* 0xe9e9 */
            {8'h00}, /* 0xe9e8 */
            {8'h00}, /* 0xe9e7 */
            {8'h00}, /* 0xe9e6 */
            {8'h00}, /* 0xe9e5 */
            {8'h00}, /* 0xe9e4 */
            {8'h00}, /* 0xe9e3 */
            {8'h00}, /* 0xe9e2 */
            {8'h00}, /* 0xe9e1 */
            {8'h00}, /* 0xe9e0 */
            {8'h00}, /* 0xe9df */
            {8'h00}, /* 0xe9de */
            {8'h00}, /* 0xe9dd */
            {8'h00}, /* 0xe9dc */
            {8'h00}, /* 0xe9db */
            {8'h00}, /* 0xe9da */
            {8'h00}, /* 0xe9d9 */
            {8'h00}, /* 0xe9d8 */
            {8'h00}, /* 0xe9d7 */
            {8'h00}, /* 0xe9d6 */
            {8'h00}, /* 0xe9d5 */
            {8'h00}, /* 0xe9d4 */
            {8'h00}, /* 0xe9d3 */
            {8'h00}, /* 0xe9d2 */
            {8'h00}, /* 0xe9d1 */
            {8'h00}, /* 0xe9d0 */
            {8'h00}, /* 0xe9cf */
            {8'h00}, /* 0xe9ce */
            {8'h00}, /* 0xe9cd */
            {8'h00}, /* 0xe9cc */
            {8'h00}, /* 0xe9cb */
            {8'h00}, /* 0xe9ca */
            {8'h00}, /* 0xe9c9 */
            {8'h00}, /* 0xe9c8 */
            {8'h00}, /* 0xe9c7 */
            {8'h00}, /* 0xe9c6 */
            {8'h00}, /* 0xe9c5 */
            {8'h00}, /* 0xe9c4 */
            {8'h00}, /* 0xe9c3 */
            {8'h00}, /* 0xe9c2 */
            {8'h00}, /* 0xe9c1 */
            {8'h00}, /* 0xe9c0 */
            {8'h00}, /* 0xe9bf */
            {8'h00}, /* 0xe9be */
            {8'h00}, /* 0xe9bd */
            {8'h00}, /* 0xe9bc */
            {8'h00}, /* 0xe9bb */
            {8'h00}, /* 0xe9ba */
            {8'h00}, /* 0xe9b9 */
            {8'h00}, /* 0xe9b8 */
            {8'h00}, /* 0xe9b7 */
            {8'h00}, /* 0xe9b6 */
            {8'h00}, /* 0xe9b5 */
            {8'h00}, /* 0xe9b4 */
            {8'h00}, /* 0xe9b3 */
            {8'h00}, /* 0xe9b2 */
            {8'h00}, /* 0xe9b1 */
            {8'h00}, /* 0xe9b0 */
            {8'h00}, /* 0xe9af */
            {8'h00}, /* 0xe9ae */
            {8'h00}, /* 0xe9ad */
            {8'h00}, /* 0xe9ac */
            {8'h00}, /* 0xe9ab */
            {8'h00}, /* 0xe9aa */
            {8'h00}, /* 0xe9a9 */
            {8'h00}, /* 0xe9a8 */
            {8'h00}, /* 0xe9a7 */
            {8'h00}, /* 0xe9a6 */
            {8'h00}, /* 0xe9a5 */
            {8'h00}, /* 0xe9a4 */
            {8'h00}, /* 0xe9a3 */
            {8'h00}, /* 0xe9a2 */
            {8'h00}, /* 0xe9a1 */
            {8'h00}, /* 0xe9a0 */
            {8'h00}, /* 0xe99f */
            {8'h00}, /* 0xe99e */
            {8'h00}, /* 0xe99d */
            {8'h00}, /* 0xe99c */
            {8'h00}, /* 0xe99b */
            {8'h00}, /* 0xe99a */
            {8'h00}, /* 0xe999 */
            {8'h00}, /* 0xe998 */
            {8'h00}, /* 0xe997 */
            {8'h00}, /* 0xe996 */
            {8'h00}, /* 0xe995 */
            {8'h00}, /* 0xe994 */
            {8'h00}, /* 0xe993 */
            {8'h00}, /* 0xe992 */
            {8'h00}, /* 0xe991 */
            {8'h00}, /* 0xe990 */
            {8'h00}, /* 0xe98f */
            {8'h00}, /* 0xe98e */
            {8'h00}, /* 0xe98d */
            {8'h00}, /* 0xe98c */
            {8'h00}, /* 0xe98b */
            {8'h00}, /* 0xe98a */
            {8'h00}, /* 0xe989 */
            {8'h00}, /* 0xe988 */
            {8'h00}, /* 0xe987 */
            {8'h00}, /* 0xe986 */
            {8'h00}, /* 0xe985 */
            {8'h00}, /* 0xe984 */
            {8'h00}, /* 0xe983 */
            {8'h00}, /* 0xe982 */
            {8'h00}, /* 0xe981 */
            {8'h00}, /* 0xe980 */
            {8'h00}, /* 0xe97f */
            {8'h00}, /* 0xe97e */
            {8'h00}, /* 0xe97d */
            {8'h00}, /* 0xe97c */
            {8'h00}, /* 0xe97b */
            {8'h00}, /* 0xe97a */
            {8'h00}, /* 0xe979 */
            {8'h00}, /* 0xe978 */
            {8'h00}, /* 0xe977 */
            {8'h00}, /* 0xe976 */
            {8'h00}, /* 0xe975 */
            {8'h00}, /* 0xe974 */
            {8'h00}, /* 0xe973 */
            {8'h00}, /* 0xe972 */
            {8'h00}, /* 0xe971 */
            {8'h00}, /* 0xe970 */
            {8'h00}, /* 0xe96f */
            {8'h00}, /* 0xe96e */
            {8'h00}, /* 0xe96d */
            {8'h00}, /* 0xe96c */
            {8'h00}, /* 0xe96b */
            {8'h00}, /* 0xe96a */
            {8'h00}, /* 0xe969 */
            {8'h00}, /* 0xe968 */
            {8'h00}, /* 0xe967 */
            {8'h00}, /* 0xe966 */
            {8'h00}, /* 0xe965 */
            {8'h00}, /* 0xe964 */
            {8'h00}, /* 0xe963 */
            {8'h00}, /* 0xe962 */
            {8'h00}, /* 0xe961 */
            {8'h00}, /* 0xe960 */
            {8'h00}, /* 0xe95f */
            {8'h00}, /* 0xe95e */
            {8'h00}, /* 0xe95d */
            {8'h00}, /* 0xe95c */
            {8'h00}, /* 0xe95b */
            {8'h00}, /* 0xe95a */
            {8'h00}, /* 0xe959 */
            {8'h00}, /* 0xe958 */
            {8'h00}, /* 0xe957 */
            {8'h00}, /* 0xe956 */
            {8'h00}, /* 0xe955 */
            {8'h00}, /* 0xe954 */
            {8'h00}, /* 0xe953 */
            {8'h00}, /* 0xe952 */
            {8'h00}, /* 0xe951 */
            {8'h00}, /* 0xe950 */
            {8'h00}, /* 0xe94f */
            {8'h00}, /* 0xe94e */
            {8'h00}, /* 0xe94d */
            {8'h00}, /* 0xe94c */
            {8'h00}, /* 0xe94b */
            {8'h00}, /* 0xe94a */
            {8'h00}, /* 0xe949 */
            {8'h00}, /* 0xe948 */
            {8'h00}, /* 0xe947 */
            {8'h00}, /* 0xe946 */
            {8'h00}, /* 0xe945 */
            {8'h00}, /* 0xe944 */
            {8'h00}, /* 0xe943 */
            {8'h00}, /* 0xe942 */
            {8'h00}, /* 0xe941 */
            {8'h00}, /* 0xe940 */
            {8'h00}, /* 0xe93f */
            {8'h00}, /* 0xe93e */
            {8'h00}, /* 0xe93d */
            {8'h00}, /* 0xe93c */
            {8'h00}, /* 0xe93b */
            {8'h00}, /* 0xe93a */
            {8'h00}, /* 0xe939 */
            {8'h00}, /* 0xe938 */
            {8'h00}, /* 0xe937 */
            {8'h00}, /* 0xe936 */
            {8'h00}, /* 0xe935 */
            {8'h00}, /* 0xe934 */
            {8'h00}, /* 0xe933 */
            {8'h00}, /* 0xe932 */
            {8'h00}, /* 0xe931 */
            {8'h00}, /* 0xe930 */
            {8'h00}, /* 0xe92f */
            {8'h00}, /* 0xe92e */
            {8'h00}, /* 0xe92d */
            {8'h00}, /* 0xe92c */
            {8'h00}, /* 0xe92b */
            {8'h00}, /* 0xe92a */
            {8'h00}, /* 0xe929 */
            {8'h00}, /* 0xe928 */
            {8'h00}, /* 0xe927 */
            {8'h00}, /* 0xe926 */
            {8'h00}, /* 0xe925 */
            {8'h00}, /* 0xe924 */
            {8'h00}, /* 0xe923 */
            {8'h00}, /* 0xe922 */
            {8'h00}, /* 0xe921 */
            {8'h00}, /* 0xe920 */
            {8'h00}, /* 0xe91f */
            {8'h00}, /* 0xe91e */
            {8'h00}, /* 0xe91d */
            {8'h00}, /* 0xe91c */
            {8'h00}, /* 0xe91b */
            {8'h00}, /* 0xe91a */
            {8'h00}, /* 0xe919 */
            {8'h00}, /* 0xe918 */
            {8'h00}, /* 0xe917 */
            {8'h00}, /* 0xe916 */
            {8'h00}, /* 0xe915 */
            {8'h00}, /* 0xe914 */
            {8'h00}, /* 0xe913 */
            {8'h00}, /* 0xe912 */
            {8'h00}, /* 0xe911 */
            {8'h00}, /* 0xe910 */
            {8'h00}, /* 0xe90f */
            {8'h00}, /* 0xe90e */
            {8'h00}, /* 0xe90d */
            {8'h00}, /* 0xe90c */
            {8'h00}, /* 0xe90b */
            {8'h00}, /* 0xe90a */
            {8'h00}, /* 0xe909 */
            {8'h00}, /* 0xe908 */
            {8'h00}, /* 0xe907 */
            {8'h00}, /* 0xe906 */
            {8'h00}, /* 0xe905 */
            {8'h00}, /* 0xe904 */
            {8'h00}, /* 0xe903 */
            {8'h00}, /* 0xe902 */
            {8'h00}, /* 0xe901 */
            {8'h00}, /* 0xe900 */
            {8'h00}, /* 0xe8ff */
            {8'h00}, /* 0xe8fe */
            {8'h00}, /* 0xe8fd */
            {8'h00}, /* 0xe8fc */
            {8'h00}, /* 0xe8fb */
            {8'h00}, /* 0xe8fa */
            {8'h00}, /* 0xe8f9 */
            {8'h00}, /* 0xe8f8 */
            {8'h00}, /* 0xe8f7 */
            {8'h00}, /* 0xe8f6 */
            {8'h00}, /* 0xe8f5 */
            {8'h00}, /* 0xe8f4 */
            {8'h00}, /* 0xe8f3 */
            {8'h00}, /* 0xe8f2 */
            {8'h00}, /* 0xe8f1 */
            {8'h00}, /* 0xe8f0 */
            {8'h00}, /* 0xe8ef */
            {8'h00}, /* 0xe8ee */
            {8'h00}, /* 0xe8ed */
            {8'h00}, /* 0xe8ec */
            {8'h00}, /* 0xe8eb */
            {8'h00}, /* 0xe8ea */
            {8'h00}, /* 0xe8e9 */
            {8'h00}, /* 0xe8e8 */
            {8'h00}, /* 0xe8e7 */
            {8'h00}, /* 0xe8e6 */
            {8'h00}, /* 0xe8e5 */
            {8'h00}, /* 0xe8e4 */
            {8'h00}, /* 0xe8e3 */
            {8'h00}, /* 0xe8e2 */
            {8'h00}, /* 0xe8e1 */
            {8'h00}, /* 0xe8e0 */
            {8'h00}, /* 0xe8df */
            {8'h00}, /* 0xe8de */
            {8'h00}, /* 0xe8dd */
            {8'h00}, /* 0xe8dc */
            {8'h00}, /* 0xe8db */
            {8'h00}, /* 0xe8da */
            {8'h00}, /* 0xe8d9 */
            {8'h00}, /* 0xe8d8 */
            {8'h00}, /* 0xe8d7 */
            {8'h00}, /* 0xe8d6 */
            {8'h00}, /* 0xe8d5 */
            {8'h00}, /* 0xe8d4 */
            {8'h00}, /* 0xe8d3 */
            {8'h00}, /* 0xe8d2 */
            {8'h00}, /* 0xe8d1 */
            {8'h00}, /* 0xe8d0 */
            {8'h00}, /* 0xe8cf */
            {8'h00}, /* 0xe8ce */
            {8'h00}, /* 0xe8cd */
            {8'h00}, /* 0xe8cc */
            {8'h00}, /* 0xe8cb */
            {8'h00}, /* 0xe8ca */
            {8'h00}, /* 0xe8c9 */
            {8'h00}, /* 0xe8c8 */
            {8'h00}, /* 0xe8c7 */
            {8'h00}, /* 0xe8c6 */
            {8'h00}, /* 0xe8c5 */
            {8'h00}, /* 0xe8c4 */
            {8'h00}, /* 0xe8c3 */
            {8'h00}, /* 0xe8c2 */
            {8'h00}, /* 0xe8c1 */
            {8'h00}, /* 0xe8c0 */
            {8'h00}, /* 0xe8bf */
            {8'h00}, /* 0xe8be */
            {8'h00}, /* 0xe8bd */
            {8'h00}, /* 0xe8bc */
            {8'h00}, /* 0xe8bb */
            {8'h00}, /* 0xe8ba */
            {8'h00}, /* 0xe8b9 */
            {8'h00}, /* 0xe8b8 */
            {8'h00}, /* 0xe8b7 */
            {8'h00}, /* 0xe8b6 */
            {8'h00}, /* 0xe8b5 */
            {8'h00}, /* 0xe8b4 */
            {8'h00}, /* 0xe8b3 */
            {8'h00}, /* 0xe8b2 */
            {8'h00}, /* 0xe8b1 */
            {8'h00}, /* 0xe8b0 */
            {8'h00}, /* 0xe8af */
            {8'h00}, /* 0xe8ae */
            {8'h00}, /* 0xe8ad */
            {8'h00}, /* 0xe8ac */
            {8'h00}, /* 0xe8ab */
            {8'h00}, /* 0xe8aa */
            {8'h00}, /* 0xe8a9 */
            {8'h00}, /* 0xe8a8 */
            {8'h00}, /* 0xe8a7 */
            {8'h00}, /* 0xe8a6 */
            {8'h00}, /* 0xe8a5 */
            {8'h00}, /* 0xe8a4 */
            {8'h00}, /* 0xe8a3 */
            {8'h00}, /* 0xe8a2 */
            {8'h00}, /* 0xe8a1 */
            {8'h00}, /* 0xe8a0 */
            {8'h00}, /* 0xe89f */
            {8'h00}, /* 0xe89e */
            {8'h00}, /* 0xe89d */
            {8'h00}, /* 0xe89c */
            {8'h00}, /* 0xe89b */
            {8'h00}, /* 0xe89a */
            {8'h00}, /* 0xe899 */
            {8'h00}, /* 0xe898 */
            {8'h00}, /* 0xe897 */
            {8'h00}, /* 0xe896 */
            {8'h00}, /* 0xe895 */
            {8'h00}, /* 0xe894 */
            {8'h00}, /* 0xe893 */
            {8'h00}, /* 0xe892 */
            {8'h00}, /* 0xe891 */
            {8'h00}, /* 0xe890 */
            {8'h00}, /* 0xe88f */
            {8'h00}, /* 0xe88e */
            {8'h00}, /* 0xe88d */
            {8'h00}, /* 0xe88c */
            {8'h00}, /* 0xe88b */
            {8'h00}, /* 0xe88a */
            {8'h00}, /* 0xe889 */
            {8'h00}, /* 0xe888 */
            {8'h00}, /* 0xe887 */
            {8'h00}, /* 0xe886 */
            {8'h00}, /* 0xe885 */
            {8'h00}, /* 0xe884 */
            {8'h00}, /* 0xe883 */
            {8'h00}, /* 0xe882 */
            {8'h00}, /* 0xe881 */
            {8'h00}, /* 0xe880 */
            {8'h00}, /* 0xe87f */
            {8'h00}, /* 0xe87e */
            {8'h00}, /* 0xe87d */
            {8'h00}, /* 0xe87c */
            {8'h00}, /* 0xe87b */
            {8'h00}, /* 0xe87a */
            {8'h00}, /* 0xe879 */
            {8'h00}, /* 0xe878 */
            {8'h00}, /* 0xe877 */
            {8'h00}, /* 0xe876 */
            {8'h00}, /* 0xe875 */
            {8'h00}, /* 0xe874 */
            {8'h00}, /* 0xe873 */
            {8'h00}, /* 0xe872 */
            {8'h00}, /* 0xe871 */
            {8'h00}, /* 0xe870 */
            {8'h00}, /* 0xe86f */
            {8'h00}, /* 0xe86e */
            {8'h00}, /* 0xe86d */
            {8'h00}, /* 0xe86c */
            {8'h00}, /* 0xe86b */
            {8'h00}, /* 0xe86a */
            {8'h00}, /* 0xe869 */
            {8'h00}, /* 0xe868 */
            {8'h00}, /* 0xe867 */
            {8'h00}, /* 0xe866 */
            {8'h00}, /* 0xe865 */
            {8'h00}, /* 0xe864 */
            {8'h00}, /* 0xe863 */
            {8'h00}, /* 0xe862 */
            {8'h00}, /* 0xe861 */
            {8'h00}, /* 0xe860 */
            {8'h00}, /* 0xe85f */
            {8'h00}, /* 0xe85e */
            {8'h00}, /* 0xe85d */
            {8'h00}, /* 0xe85c */
            {8'h00}, /* 0xe85b */
            {8'h00}, /* 0xe85a */
            {8'h00}, /* 0xe859 */
            {8'h00}, /* 0xe858 */
            {8'h00}, /* 0xe857 */
            {8'h00}, /* 0xe856 */
            {8'h00}, /* 0xe855 */
            {8'h00}, /* 0xe854 */
            {8'h00}, /* 0xe853 */
            {8'h00}, /* 0xe852 */
            {8'h00}, /* 0xe851 */
            {8'h00}, /* 0xe850 */
            {8'h00}, /* 0xe84f */
            {8'h00}, /* 0xe84e */
            {8'h00}, /* 0xe84d */
            {8'h00}, /* 0xe84c */
            {8'h00}, /* 0xe84b */
            {8'h00}, /* 0xe84a */
            {8'h00}, /* 0xe849 */
            {8'h00}, /* 0xe848 */
            {8'h00}, /* 0xe847 */
            {8'h00}, /* 0xe846 */
            {8'h00}, /* 0xe845 */
            {8'h00}, /* 0xe844 */
            {8'h00}, /* 0xe843 */
            {8'h00}, /* 0xe842 */
            {8'h00}, /* 0xe841 */
            {8'h00}, /* 0xe840 */
            {8'h00}, /* 0xe83f */
            {8'h00}, /* 0xe83e */
            {8'h00}, /* 0xe83d */
            {8'h00}, /* 0xe83c */
            {8'h00}, /* 0xe83b */
            {8'h00}, /* 0xe83a */
            {8'h00}, /* 0xe839 */
            {8'h00}, /* 0xe838 */
            {8'h00}, /* 0xe837 */
            {8'h00}, /* 0xe836 */
            {8'h00}, /* 0xe835 */
            {8'h00}, /* 0xe834 */
            {8'h00}, /* 0xe833 */
            {8'h00}, /* 0xe832 */
            {8'h00}, /* 0xe831 */
            {8'h00}, /* 0xe830 */
            {8'h00}, /* 0xe82f */
            {8'h00}, /* 0xe82e */
            {8'h00}, /* 0xe82d */
            {8'h00}, /* 0xe82c */
            {8'h00}, /* 0xe82b */
            {8'h00}, /* 0xe82a */
            {8'h00}, /* 0xe829 */
            {8'h00}, /* 0xe828 */
            {8'h00}, /* 0xe827 */
            {8'h00}, /* 0xe826 */
            {8'h00}, /* 0xe825 */
            {8'h00}, /* 0xe824 */
            {8'h00}, /* 0xe823 */
            {8'h00}, /* 0xe822 */
            {8'h00}, /* 0xe821 */
            {8'h00}, /* 0xe820 */
            {8'h00}, /* 0xe81f */
            {8'h00}, /* 0xe81e */
            {8'h00}, /* 0xe81d */
            {8'h00}, /* 0xe81c */
            {8'h00}, /* 0xe81b */
            {8'h00}, /* 0xe81a */
            {8'h00}, /* 0xe819 */
            {8'h00}, /* 0xe818 */
            {8'h00}, /* 0xe817 */
            {8'h00}, /* 0xe816 */
            {8'h00}, /* 0xe815 */
            {8'h00}, /* 0xe814 */
            {8'h00}, /* 0xe813 */
            {8'h00}, /* 0xe812 */
            {8'h00}, /* 0xe811 */
            {8'h00}, /* 0xe810 */
            {8'h00}, /* 0xe80f */
            {8'h00}, /* 0xe80e */
            {8'h00}, /* 0xe80d */
            {8'h00}, /* 0xe80c */
            {8'h00}, /* 0xe80b */
            {8'h00}, /* 0xe80a */
            {8'h00}, /* 0xe809 */
            {8'h00}, /* 0xe808 */
            {8'h00}, /* 0xe807 */
            {8'h00}, /* 0xe806 */
            {8'h00}, /* 0xe805 */
            {8'h00}, /* 0xe804 */
            {8'h00}, /* 0xe803 */
            {8'h00}, /* 0xe802 */
            {8'h00}, /* 0xe801 */
            {8'h00}, /* 0xe800 */
            {8'h00}, /* 0xe7ff */
            {8'h00}, /* 0xe7fe */
            {8'h00}, /* 0xe7fd */
            {8'h00}, /* 0xe7fc */
            {8'h00}, /* 0xe7fb */
            {8'h00}, /* 0xe7fa */
            {8'h00}, /* 0xe7f9 */
            {8'h00}, /* 0xe7f8 */
            {8'h00}, /* 0xe7f7 */
            {8'h00}, /* 0xe7f6 */
            {8'h00}, /* 0xe7f5 */
            {8'h00}, /* 0xe7f4 */
            {8'h00}, /* 0xe7f3 */
            {8'h00}, /* 0xe7f2 */
            {8'h00}, /* 0xe7f1 */
            {8'h00}, /* 0xe7f0 */
            {8'h00}, /* 0xe7ef */
            {8'h00}, /* 0xe7ee */
            {8'h00}, /* 0xe7ed */
            {8'h00}, /* 0xe7ec */
            {8'h00}, /* 0xe7eb */
            {8'h00}, /* 0xe7ea */
            {8'h00}, /* 0xe7e9 */
            {8'h00}, /* 0xe7e8 */
            {8'h00}, /* 0xe7e7 */
            {8'h00}, /* 0xe7e6 */
            {8'h00}, /* 0xe7e5 */
            {8'h00}, /* 0xe7e4 */
            {8'h00}, /* 0xe7e3 */
            {8'h00}, /* 0xe7e2 */
            {8'h00}, /* 0xe7e1 */
            {8'h00}, /* 0xe7e0 */
            {8'h00}, /* 0xe7df */
            {8'h00}, /* 0xe7de */
            {8'h00}, /* 0xe7dd */
            {8'h00}, /* 0xe7dc */
            {8'h00}, /* 0xe7db */
            {8'h00}, /* 0xe7da */
            {8'h00}, /* 0xe7d9 */
            {8'h00}, /* 0xe7d8 */
            {8'h00}, /* 0xe7d7 */
            {8'h00}, /* 0xe7d6 */
            {8'h00}, /* 0xe7d5 */
            {8'h00}, /* 0xe7d4 */
            {8'h00}, /* 0xe7d3 */
            {8'h00}, /* 0xe7d2 */
            {8'h00}, /* 0xe7d1 */
            {8'h00}, /* 0xe7d0 */
            {8'h00}, /* 0xe7cf */
            {8'h00}, /* 0xe7ce */
            {8'h00}, /* 0xe7cd */
            {8'h00}, /* 0xe7cc */
            {8'h00}, /* 0xe7cb */
            {8'h00}, /* 0xe7ca */
            {8'h00}, /* 0xe7c9 */
            {8'h00}, /* 0xe7c8 */
            {8'h00}, /* 0xe7c7 */
            {8'h00}, /* 0xe7c6 */
            {8'h00}, /* 0xe7c5 */
            {8'h00}, /* 0xe7c4 */
            {8'h00}, /* 0xe7c3 */
            {8'h00}, /* 0xe7c2 */
            {8'h00}, /* 0xe7c1 */
            {8'h00}, /* 0xe7c0 */
            {8'h00}, /* 0xe7bf */
            {8'h00}, /* 0xe7be */
            {8'h00}, /* 0xe7bd */
            {8'h00}, /* 0xe7bc */
            {8'h00}, /* 0xe7bb */
            {8'h00}, /* 0xe7ba */
            {8'h00}, /* 0xe7b9 */
            {8'h00}, /* 0xe7b8 */
            {8'h00}, /* 0xe7b7 */
            {8'h00}, /* 0xe7b6 */
            {8'h00}, /* 0xe7b5 */
            {8'h00}, /* 0xe7b4 */
            {8'h00}, /* 0xe7b3 */
            {8'h00}, /* 0xe7b2 */
            {8'h00}, /* 0xe7b1 */
            {8'h00}, /* 0xe7b0 */
            {8'h00}, /* 0xe7af */
            {8'h00}, /* 0xe7ae */
            {8'h00}, /* 0xe7ad */
            {8'h00}, /* 0xe7ac */
            {8'h00}, /* 0xe7ab */
            {8'h00}, /* 0xe7aa */
            {8'h00}, /* 0xe7a9 */
            {8'h00}, /* 0xe7a8 */
            {8'h00}, /* 0xe7a7 */
            {8'h00}, /* 0xe7a6 */
            {8'h00}, /* 0xe7a5 */
            {8'h00}, /* 0xe7a4 */
            {8'h00}, /* 0xe7a3 */
            {8'h00}, /* 0xe7a2 */
            {8'h00}, /* 0xe7a1 */
            {8'h00}, /* 0xe7a0 */
            {8'h00}, /* 0xe79f */
            {8'h00}, /* 0xe79e */
            {8'h00}, /* 0xe79d */
            {8'h00}, /* 0xe79c */
            {8'h00}, /* 0xe79b */
            {8'h00}, /* 0xe79a */
            {8'h00}, /* 0xe799 */
            {8'h00}, /* 0xe798 */
            {8'h00}, /* 0xe797 */
            {8'h00}, /* 0xe796 */
            {8'h00}, /* 0xe795 */
            {8'h00}, /* 0xe794 */
            {8'h00}, /* 0xe793 */
            {8'h00}, /* 0xe792 */
            {8'h00}, /* 0xe791 */
            {8'h00}, /* 0xe790 */
            {8'h00}, /* 0xe78f */
            {8'h00}, /* 0xe78e */
            {8'h00}, /* 0xe78d */
            {8'h00}, /* 0xe78c */
            {8'h00}, /* 0xe78b */
            {8'h00}, /* 0xe78a */
            {8'h00}, /* 0xe789 */
            {8'h00}, /* 0xe788 */
            {8'h00}, /* 0xe787 */
            {8'h00}, /* 0xe786 */
            {8'h00}, /* 0xe785 */
            {8'h00}, /* 0xe784 */
            {8'h00}, /* 0xe783 */
            {8'h00}, /* 0xe782 */
            {8'h00}, /* 0xe781 */
            {8'h00}, /* 0xe780 */
            {8'h00}, /* 0xe77f */
            {8'h00}, /* 0xe77e */
            {8'h00}, /* 0xe77d */
            {8'h00}, /* 0xe77c */
            {8'h00}, /* 0xe77b */
            {8'h00}, /* 0xe77a */
            {8'h00}, /* 0xe779 */
            {8'h00}, /* 0xe778 */
            {8'h00}, /* 0xe777 */
            {8'h00}, /* 0xe776 */
            {8'h00}, /* 0xe775 */
            {8'h00}, /* 0xe774 */
            {8'h00}, /* 0xe773 */
            {8'h00}, /* 0xe772 */
            {8'h00}, /* 0xe771 */
            {8'h00}, /* 0xe770 */
            {8'h00}, /* 0xe76f */
            {8'h00}, /* 0xe76e */
            {8'h00}, /* 0xe76d */
            {8'h00}, /* 0xe76c */
            {8'h00}, /* 0xe76b */
            {8'h00}, /* 0xe76a */
            {8'h00}, /* 0xe769 */
            {8'h00}, /* 0xe768 */
            {8'h00}, /* 0xe767 */
            {8'h00}, /* 0xe766 */
            {8'h00}, /* 0xe765 */
            {8'h00}, /* 0xe764 */
            {8'h00}, /* 0xe763 */
            {8'h00}, /* 0xe762 */
            {8'h00}, /* 0xe761 */
            {8'h00}, /* 0xe760 */
            {8'h00}, /* 0xe75f */
            {8'h00}, /* 0xe75e */
            {8'h00}, /* 0xe75d */
            {8'h00}, /* 0xe75c */
            {8'h00}, /* 0xe75b */
            {8'h00}, /* 0xe75a */
            {8'h00}, /* 0xe759 */
            {8'h00}, /* 0xe758 */
            {8'h00}, /* 0xe757 */
            {8'h00}, /* 0xe756 */
            {8'h00}, /* 0xe755 */
            {8'h00}, /* 0xe754 */
            {8'h00}, /* 0xe753 */
            {8'h00}, /* 0xe752 */
            {8'h00}, /* 0xe751 */
            {8'h00}, /* 0xe750 */
            {8'h00}, /* 0xe74f */
            {8'h00}, /* 0xe74e */
            {8'h00}, /* 0xe74d */
            {8'h00}, /* 0xe74c */
            {8'h00}, /* 0xe74b */
            {8'h00}, /* 0xe74a */
            {8'h00}, /* 0xe749 */
            {8'h00}, /* 0xe748 */
            {8'h00}, /* 0xe747 */
            {8'h00}, /* 0xe746 */
            {8'h00}, /* 0xe745 */
            {8'h00}, /* 0xe744 */
            {8'h00}, /* 0xe743 */
            {8'h00}, /* 0xe742 */
            {8'h00}, /* 0xe741 */
            {8'h00}, /* 0xe740 */
            {8'h00}, /* 0xe73f */
            {8'h00}, /* 0xe73e */
            {8'h00}, /* 0xe73d */
            {8'h00}, /* 0xe73c */
            {8'h00}, /* 0xe73b */
            {8'h00}, /* 0xe73a */
            {8'h00}, /* 0xe739 */
            {8'h00}, /* 0xe738 */
            {8'h00}, /* 0xe737 */
            {8'h00}, /* 0xe736 */
            {8'h00}, /* 0xe735 */
            {8'h00}, /* 0xe734 */
            {8'h00}, /* 0xe733 */
            {8'h00}, /* 0xe732 */
            {8'h00}, /* 0xe731 */
            {8'h00}, /* 0xe730 */
            {8'h00}, /* 0xe72f */
            {8'h00}, /* 0xe72e */
            {8'h00}, /* 0xe72d */
            {8'h00}, /* 0xe72c */
            {8'h00}, /* 0xe72b */
            {8'h00}, /* 0xe72a */
            {8'h00}, /* 0xe729 */
            {8'h00}, /* 0xe728 */
            {8'h00}, /* 0xe727 */
            {8'h00}, /* 0xe726 */
            {8'h00}, /* 0xe725 */
            {8'h00}, /* 0xe724 */
            {8'h00}, /* 0xe723 */
            {8'h00}, /* 0xe722 */
            {8'h00}, /* 0xe721 */
            {8'h00}, /* 0xe720 */
            {8'h00}, /* 0xe71f */
            {8'h00}, /* 0xe71e */
            {8'h00}, /* 0xe71d */
            {8'h00}, /* 0xe71c */
            {8'h00}, /* 0xe71b */
            {8'h00}, /* 0xe71a */
            {8'h00}, /* 0xe719 */
            {8'h00}, /* 0xe718 */
            {8'h00}, /* 0xe717 */
            {8'h00}, /* 0xe716 */
            {8'h00}, /* 0xe715 */
            {8'h00}, /* 0xe714 */
            {8'h00}, /* 0xe713 */
            {8'h00}, /* 0xe712 */
            {8'h00}, /* 0xe711 */
            {8'h00}, /* 0xe710 */
            {8'h00}, /* 0xe70f */
            {8'h00}, /* 0xe70e */
            {8'h00}, /* 0xe70d */
            {8'h00}, /* 0xe70c */
            {8'h00}, /* 0xe70b */
            {8'h00}, /* 0xe70a */
            {8'h00}, /* 0xe709 */
            {8'h00}, /* 0xe708 */
            {8'h00}, /* 0xe707 */
            {8'h00}, /* 0xe706 */
            {8'h00}, /* 0xe705 */
            {8'h00}, /* 0xe704 */
            {8'h00}, /* 0xe703 */
            {8'h00}, /* 0xe702 */
            {8'h00}, /* 0xe701 */
            {8'h00}, /* 0xe700 */
            {8'h00}, /* 0xe6ff */
            {8'h00}, /* 0xe6fe */
            {8'h00}, /* 0xe6fd */
            {8'h00}, /* 0xe6fc */
            {8'h00}, /* 0xe6fb */
            {8'h00}, /* 0xe6fa */
            {8'h00}, /* 0xe6f9 */
            {8'h00}, /* 0xe6f8 */
            {8'h00}, /* 0xe6f7 */
            {8'h00}, /* 0xe6f6 */
            {8'h00}, /* 0xe6f5 */
            {8'h00}, /* 0xe6f4 */
            {8'h00}, /* 0xe6f3 */
            {8'h00}, /* 0xe6f2 */
            {8'h00}, /* 0xe6f1 */
            {8'h00}, /* 0xe6f0 */
            {8'h00}, /* 0xe6ef */
            {8'h00}, /* 0xe6ee */
            {8'h00}, /* 0xe6ed */
            {8'h00}, /* 0xe6ec */
            {8'h00}, /* 0xe6eb */
            {8'h00}, /* 0xe6ea */
            {8'h00}, /* 0xe6e9 */
            {8'h00}, /* 0xe6e8 */
            {8'h00}, /* 0xe6e7 */
            {8'h00}, /* 0xe6e6 */
            {8'h00}, /* 0xe6e5 */
            {8'h00}, /* 0xe6e4 */
            {8'h00}, /* 0xe6e3 */
            {8'h00}, /* 0xe6e2 */
            {8'h00}, /* 0xe6e1 */
            {8'h00}, /* 0xe6e0 */
            {8'h00}, /* 0xe6df */
            {8'h00}, /* 0xe6de */
            {8'h00}, /* 0xe6dd */
            {8'h00}, /* 0xe6dc */
            {8'h00}, /* 0xe6db */
            {8'h00}, /* 0xe6da */
            {8'h00}, /* 0xe6d9 */
            {8'h00}, /* 0xe6d8 */
            {8'h00}, /* 0xe6d7 */
            {8'h00}, /* 0xe6d6 */
            {8'h00}, /* 0xe6d5 */
            {8'h00}, /* 0xe6d4 */
            {8'h00}, /* 0xe6d3 */
            {8'h00}, /* 0xe6d2 */
            {8'h00}, /* 0xe6d1 */
            {8'h00}, /* 0xe6d0 */
            {8'h00}, /* 0xe6cf */
            {8'h00}, /* 0xe6ce */
            {8'h00}, /* 0xe6cd */
            {8'h00}, /* 0xe6cc */
            {8'h00}, /* 0xe6cb */
            {8'h00}, /* 0xe6ca */
            {8'h00}, /* 0xe6c9 */
            {8'h00}, /* 0xe6c8 */
            {8'h00}, /* 0xe6c7 */
            {8'h00}, /* 0xe6c6 */
            {8'h00}, /* 0xe6c5 */
            {8'h00}, /* 0xe6c4 */
            {8'h00}, /* 0xe6c3 */
            {8'h00}, /* 0xe6c2 */
            {8'h00}, /* 0xe6c1 */
            {8'h00}, /* 0xe6c0 */
            {8'h00}, /* 0xe6bf */
            {8'h00}, /* 0xe6be */
            {8'h00}, /* 0xe6bd */
            {8'h00}, /* 0xe6bc */
            {8'h00}, /* 0xe6bb */
            {8'h00}, /* 0xe6ba */
            {8'h00}, /* 0xe6b9 */
            {8'h00}, /* 0xe6b8 */
            {8'h00}, /* 0xe6b7 */
            {8'h00}, /* 0xe6b6 */
            {8'h00}, /* 0xe6b5 */
            {8'h00}, /* 0xe6b4 */
            {8'h00}, /* 0xe6b3 */
            {8'h00}, /* 0xe6b2 */
            {8'h00}, /* 0xe6b1 */
            {8'h00}, /* 0xe6b0 */
            {8'h00}, /* 0xe6af */
            {8'h00}, /* 0xe6ae */
            {8'h00}, /* 0xe6ad */
            {8'h00}, /* 0xe6ac */
            {8'h00}, /* 0xe6ab */
            {8'h00}, /* 0xe6aa */
            {8'h00}, /* 0xe6a9 */
            {8'h00}, /* 0xe6a8 */
            {8'h00}, /* 0xe6a7 */
            {8'h00}, /* 0xe6a6 */
            {8'h00}, /* 0xe6a5 */
            {8'h00}, /* 0xe6a4 */
            {8'h00}, /* 0xe6a3 */
            {8'h00}, /* 0xe6a2 */
            {8'h00}, /* 0xe6a1 */
            {8'h00}, /* 0xe6a0 */
            {8'h00}, /* 0xe69f */
            {8'h00}, /* 0xe69e */
            {8'h00}, /* 0xe69d */
            {8'h00}, /* 0xe69c */
            {8'h00}, /* 0xe69b */
            {8'h00}, /* 0xe69a */
            {8'h00}, /* 0xe699 */
            {8'h00}, /* 0xe698 */
            {8'h00}, /* 0xe697 */
            {8'h00}, /* 0xe696 */
            {8'h00}, /* 0xe695 */
            {8'h00}, /* 0xe694 */
            {8'h00}, /* 0xe693 */
            {8'h00}, /* 0xe692 */
            {8'h00}, /* 0xe691 */
            {8'h00}, /* 0xe690 */
            {8'h00}, /* 0xe68f */
            {8'h00}, /* 0xe68e */
            {8'h00}, /* 0xe68d */
            {8'h00}, /* 0xe68c */
            {8'h00}, /* 0xe68b */
            {8'h00}, /* 0xe68a */
            {8'h00}, /* 0xe689 */
            {8'h00}, /* 0xe688 */
            {8'h00}, /* 0xe687 */
            {8'h00}, /* 0xe686 */
            {8'h00}, /* 0xe685 */
            {8'h00}, /* 0xe684 */
            {8'h00}, /* 0xe683 */
            {8'h00}, /* 0xe682 */
            {8'h00}, /* 0xe681 */
            {8'h00}, /* 0xe680 */
            {8'h00}, /* 0xe67f */
            {8'h00}, /* 0xe67e */
            {8'h00}, /* 0xe67d */
            {8'h00}, /* 0xe67c */
            {8'h00}, /* 0xe67b */
            {8'h00}, /* 0xe67a */
            {8'h00}, /* 0xe679 */
            {8'h00}, /* 0xe678 */
            {8'h00}, /* 0xe677 */
            {8'h00}, /* 0xe676 */
            {8'h00}, /* 0xe675 */
            {8'h00}, /* 0xe674 */
            {8'h00}, /* 0xe673 */
            {8'h00}, /* 0xe672 */
            {8'h00}, /* 0xe671 */
            {8'h00}, /* 0xe670 */
            {8'h00}, /* 0xe66f */
            {8'h00}, /* 0xe66e */
            {8'h00}, /* 0xe66d */
            {8'h00}, /* 0xe66c */
            {8'h00}, /* 0xe66b */
            {8'h00}, /* 0xe66a */
            {8'h00}, /* 0xe669 */
            {8'h00}, /* 0xe668 */
            {8'h00}, /* 0xe667 */
            {8'h00}, /* 0xe666 */
            {8'h00}, /* 0xe665 */
            {8'h00}, /* 0xe664 */
            {8'h00}, /* 0xe663 */
            {8'h00}, /* 0xe662 */
            {8'h00}, /* 0xe661 */
            {8'h00}, /* 0xe660 */
            {8'h00}, /* 0xe65f */
            {8'h00}, /* 0xe65e */
            {8'h00}, /* 0xe65d */
            {8'h00}, /* 0xe65c */
            {8'h00}, /* 0xe65b */
            {8'h00}, /* 0xe65a */
            {8'h00}, /* 0xe659 */
            {8'h00}, /* 0xe658 */
            {8'h00}, /* 0xe657 */
            {8'h00}, /* 0xe656 */
            {8'h00}, /* 0xe655 */
            {8'h00}, /* 0xe654 */
            {8'h00}, /* 0xe653 */
            {8'h00}, /* 0xe652 */
            {8'h00}, /* 0xe651 */
            {8'h00}, /* 0xe650 */
            {8'h00}, /* 0xe64f */
            {8'h00}, /* 0xe64e */
            {8'h00}, /* 0xe64d */
            {8'h00}, /* 0xe64c */
            {8'h00}, /* 0xe64b */
            {8'h00}, /* 0xe64a */
            {8'h00}, /* 0xe649 */
            {8'h00}, /* 0xe648 */
            {8'h00}, /* 0xe647 */
            {8'h00}, /* 0xe646 */
            {8'h00}, /* 0xe645 */
            {8'h00}, /* 0xe644 */
            {8'h00}, /* 0xe643 */
            {8'h00}, /* 0xe642 */
            {8'h00}, /* 0xe641 */
            {8'h00}, /* 0xe640 */
            {8'h00}, /* 0xe63f */
            {8'h00}, /* 0xe63e */
            {8'h00}, /* 0xe63d */
            {8'h00}, /* 0xe63c */
            {8'h00}, /* 0xe63b */
            {8'h00}, /* 0xe63a */
            {8'h00}, /* 0xe639 */
            {8'h00}, /* 0xe638 */
            {8'h00}, /* 0xe637 */
            {8'h00}, /* 0xe636 */
            {8'h00}, /* 0xe635 */
            {8'h00}, /* 0xe634 */
            {8'h00}, /* 0xe633 */
            {8'h00}, /* 0xe632 */
            {8'h00}, /* 0xe631 */
            {8'h00}, /* 0xe630 */
            {8'h00}, /* 0xe62f */
            {8'h00}, /* 0xe62e */
            {8'h00}, /* 0xe62d */
            {8'h00}, /* 0xe62c */
            {8'h00}, /* 0xe62b */
            {8'h00}, /* 0xe62a */
            {8'h00}, /* 0xe629 */
            {8'h00}, /* 0xe628 */
            {8'h00}, /* 0xe627 */
            {8'h00}, /* 0xe626 */
            {8'h00}, /* 0xe625 */
            {8'h00}, /* 0xe624 */
            {8'h00}, /* 0xe623 */
            {8'h00}, /* 0xe622 */
            {8'h00}, /* 0xe621 */
            {8'h00}, /* 0xe620 */
            {8'h00}, /* 0xe61f */
            {8'h00}, /* 0xe61e */
            {8'h00}, /* 0xe61d */
            {8'h00}, /* 0xe61c */
            {8'h00}, /* 0xe61b */
            {8'h00}, /* 0xe61a */
            {8'h00}, /* 0xe619 */
            {8'h00}, /* 0xe618 */
            {8'h00}, /* 0xe617 */
            {8'h00}, /* 0xe616 */
            {8'h00}, /* 0xe615 */
            {8'h00}, /* 0xe614 */
            {8'h00}, /* 0xe613 */
            {8'h00}, /* 0xe612 */
            {8'h00}, /* 0xe611 */
            {8'h00}, /* 0xe610 */
            {8'h00}, /* 0xe60f */
            {8'h00}, /* 0xe60e */
            {8'h00}, /* 0xe60d */
            {8'h00}, /* 0xe60c */
            {8'h00}, /* 0xe60b */
            {8'h00}, /* 0xe60a */
            {8'h00}, /* 0xe609 */
            {8'h00}, /* 0xe608 */
            {8'h00}, /* 0xe607 */
            {8'h00}, /* 0xe606 */
            {8'h00}, /* 0xe605 */
            {8'h00}, /* 0xe604 */
            {8'h00}, /* 0xe603 */
            {8'h00}, /* 0xe602 */
            {8'h00}, /* 0xe601 */
            {8'h00}, /* 0xe600 */
            {8'h00}, /* 0xe5ff */
            {8'h00}, /* 0xe5fe */
            {8'h00}, /* 0xe5fd */
            {8'h00}, /* 0xe5fc */
            {8'h00}, /* 0xe5fb */
            {8'h00}, /* 0xe5fa */
            {8'h00}, /* 0xe5f9 */
            {8'h00}, /* 0xe5f8 */
            {8'h00}, /* 0xe5f7 */
            {8'h00}, /* 0xe5f6 */
            {8'h00}, /* 0xe5f5 */
            {8'h00}, /* 0xe5f4 */
            {8'h00}, /* 0xe5f3 */
            {8'h00}, /* 0xe5f2 */
            {8'h00}, /* 0xe5f1 */
            {8'h00}, /* 0xe5f0 */
            {8'h00}, /* 0xe5ef */
            {8'h00}, /* 0xe5ee */
            {8'h00}, /* 0xe5ed */
            {8'h00}, /* 0xe5ec */
            {8'h00}, /* 0xe5eb */
            {8'h00}, /* 0xe5ea */
            {8'h00}, /* 0xe5e9 */
            {8'h00}, /* 0xe5e8 */
            {8'h00}, /* 0xe5e7 */
            {8'h00}, /* 0xe5e6 */
            {8'h00}, /* 0xe5e5 */
            {8'h00}, /* 0xe5e4 */
            {8'h00}, /* 0xe5e3 */
            {8'h00}, /* 0xe5e2 */
            {8'h00}, /* 0xe5e1 */
            {8'h00}, /* 0xe5e0 */
            {8'h00}, /* 0xe5df */
            {8'h00}, /* 0xe5de */
            {8'h00}, /* 0xe5dd */
            {8'h00}, /* 0xe5dc */
            {8'h00}, /* 0xe5db */
            {8'h00}, /* 0xe5da */
            {8'h00}, /* 0xe5d9 */
            {8'h00}, /* 0xe5d8 */
            {8'h00}, /* 0xe5d7 */
            {8'h00}, /* 0xe5d6 */
            {8'h00}, /* 0xe5d5 */
            {8'h00}, /* 0xe5d4 */
            {8'h00}, /* 0xe5d3 */
            {8'h00}, /* 0xe5d2 */
            {8'h00}, /* 0xe5d1 */
            {8'h00}, /* 0xe5d0 */
            {8'h00}, /* 0xe5cf */
            {8'h00}, /* 0xe5ce */
            {8'h00}, /* 0xe5cd */
            {8'h00}, /* 0xe5cc */
            {8'h00}, /* 0xe5cb */
            {8'h00}, /* 0xe5ca */
            {8'h00}, /* 0xe5c9 */
            {8'h00}, /* 0xe5c8 */
            {8'h00}, /* 0xe5c7 */
            {8'h00}, /* 0xe5c6 */
            {8'h00}, /* 0xe5c5 */
            {8'h00}, /* 0xe5c4 */
            {8'h00}, /* 0xe5c3 */
            {8'h00}, /* 0xe5c2 */
            {8'h00}, /* 0xe5c1 */
            {8'h00}, /* 0xe5c0 */
            {8'h00}, /* 0xe5bf */
            {8'h00}, /* 0xe5be */
            {8'h00}, /* 0xe5bd */
            {8'h00}, /* 0xe5bc */
            {8'h00}, /* 0xe5bb */
            {8'h00}, /* 0xe5ba */
            {8'h00}, /* 0xe5b9 */
            {8'h00}, /* 0xe5b8 */
            {8'h00}, /* 0xe5b7 */
            {8'h00}, /* 0xe5b6 */
            {8'h00}, /* 0xe5b5 */
            {8'h00}, /* 0xe5b4 */
            {8'h00}, /* 0xe5b3 */
            {8'h00}, /* 0xe5b2 */
            {8'h00}, /* 0xe5b1 */
            {8'h00}, /* 0xe5b0 */
            {8'h00}, /* 0xe5af */
            {8'h00}, /* 0xe5ae */
            {8'h00}, /* 0xe5ad */
            {8'h00}, /* 0xe5ac */
            {8'h00}, /* 0xe5ab */
            {8'h00}, /* 0xe5aa */
            {8'h00}, /* 0xe5a9 */
            {8'h00}, /* 0xe5a8 */
            {8'h00}, /* 0xe5a7 */
            {8'h00}, /* 0xe5a6 */
            {8'h00}, /* 0xe5a5 */
            {8'h00}, /* 0xe5a4 */
            {8'h00}, /* 0xe5a3 */
            {8'h00}, /* 0xe5a2 */
            {8'h00}, /* 0xe5a1 */
            {8'h00}, /* 0xe5a0 */
            {8'h00}, /* 0xe59f */
            {8'h00}, /* 0xe59e */
            {8'h00}, /* 0xe59d */
            {8'h00}, /* 0xe59c */
            {8'h00}, /* 0xe59b */
            {8'h00}, /* 0xe59a */
            {8'h00}, /* 0xe599 */
            {8'h00}, /* 0xe598 */
            {8'h00}, /* 0xe597 */
            {8'h00}, /* 0xe596 */
            {8'h00}, /* 0xe595 */
            {8'h00}, /* 0xe594 */
            {8'h00}, /* 0xe593 */
            {8'h00}, /* 0xe592 */
            {8'h00}, /* 0xe591 */
            {8'h00}, /* 0xe590 */
            {8'h00}, /* 0xe58f */
            {8'h00}, /* 0xe58e */
            {8'h00}, /* 0xe58d */
            {8'h00}, /* 0xe58c */
            {8'h00}, /* 0xe58b */
            {8'h00}, /* 0xe58a */
            {8'h00}, /* 0xe589 */
            {8'h00}, /* 0xe588 */
            {8'h00}, /* 0xe587 */
            {8'h00}, /* 0xe586 */
            {8'h00}, /* 0xe585 */
            {8'h00}, /* 0xe584 */
            {8'h00}, /* 0xe583 */
            {8'h00}, /* 0xe582 */
            {8'h00}, /* 0xe581 */
            {8'h00}, /* 0xe580 */
            {8'h00}, /* 0xe57f */
            {8'h00}, /* 0xe57e */
            {8'h00}, /* 0xe57d */
            {8'h00}, /* 0xe57c */
            {8'h00}, /* 0xe57b */
            {8'h00}, /* 0xe57a */
            {8'h00}, /* 0xe579 */
            {8'h00}, /* 0xe578 */
            {8'h00}, /* 0xe577 */
            {8'h00}, /* 0xe576 */
            {8'h00}, /* 0xe575 */
            {8'h00}, /* 0xe574 */
            {8'h00}, /* 0xe573 */
            {8'h00}, /* 0xe572 */
            {8'h00}, /* 0xe571 */
            {8'h00}, /* 0xe570 */
            {8'h00}, /* 0xe56f */
            {8'h00}, /* 0xe56e */
            {8'h00}, /* 0xe56d */
            {8'h00}, /* 0xe56c */
            {8'h00}, /* 0xe56b */
            {8'h00}, /* 0xe56a */
            {8'h00}, /* 0xe569 */
            {8'h00}, /* 0xe568 */
            {8'h00}, /* 0xe567 */
            {8'h00}, /* 0xe566 */
            {8'h00}, /* 0xe565 */
            {8'h00}, /* 0xe564 */
            {8'h00}, /* 0xe563 */
            {8'h00}, /* 0xe562 */
            {8'h00}, /* 0xe561 */
            {8'h00}, /* 0xe560 */
            {8'h00}, /* 0xe55f */
            {8'h00}, /* 0xe55e */
            {8'h00}, /* 0xe55d */
            {8'h00}, /* 0xe55c */
            {8'h00}, /* 0xe55b */
            {8'h00}, /* 0xe55a */
            {8'h00}, /* 0xe559 */
            {8'h00}, /* 0xe558 */
            {8'h00}, /* 0xe557 */
            {8'h00}, /* 0xe556 */
            {8'h00}, /* 0xe555 */
            {8'h00}, /* 0xe554 */
            {8'h00}, /* 0xe553 */
            {8'h00}, /* 0xe552 */
            {8'h00}, /* 0xe551 */
            {8'h00}, /* 0xe550 */
            {8'h00}, /* 0xe54f */
            {8'h00}, /* 0xe54e */
            {8'h00}, /* 0xe54d */
            {8'h00}, /* 0xe54c */
            {8'h00}, /* 0xe54b */
            {8'h00}, /* 0xe54a */
            {8'h00}, /* 0xe549 */
            {8'h00}, /* 0xe548 */
            {8'h00}, /* 0xe547 */
            {8'h00}, /* 0xe546 */
            {8'h00}, /* 0xe545 */
            {8'h00}, /* 0xe544 */
            {8'h00}, /* 0xe543 */
            {8'h00}, /* 0xe542 */
            {8'h00}, /* 0xe541 */
            {8'h00}, /* 0xe540 */
            {8'h00}, /* 0xe53f */
            {8'h00}, /* 0xe53e */
            {8'h00}, /* 0xe53d */
            {8'h00}, /* 0xe53c */
            {8'h00}, /* 0xe53b */
            {8'h00}, /* 0xe53a */
            {8'h00}, /* 0xe539 */
            {8'h00}, /* 0xe538 */
            {8'h00}, /* 0xe537 */
            {8'h00}, /* 0xe536 */
            {8'h00}, /* 0xe535 */
            {8'h00}, /* 0xe534 */
            {8'h00}, /* 0xe533 */
            {8'h00}, /* 0xe532 */
            {8'h00}, /* 0xe531 */
            {8'h00}, /* 0xe530 */
            {8'h00}, /* 0xe52f */
            {8'h00}, /* 0xe52e */
            {8'h00}, /* 0xe52d */
            {8'h00}, /* 0xe52c */
            {8'h00}, /* 0xe52b */
            {8'h00}, /* 0xe52a */
            {8'h00}, /* 0xe529 */
            {8'h00}, /* 0xe528 */
            {8'h00}, /* 0xe527 */
            {8'h00}, /* 0xe526 */
            {8'h00}, /* 0xe525 */
            {8'h00}, /* 0xe524 */
            {8'h00}, /* 0xe523 */
            {8'h00}, /* 0xe522 */
            {8'h00}, /* 0xe521 */
            {8'h00}, /* 0xe520 */
            {8'h00}, /* 0xe51f */
            {8'h00}, /* 0xe51e */
            {8'h00}, /* 0xe51d */
            {8'h00}, /* 0xe51c */
            {8'h00}, /* 0xe51b */
            {8'h00}, /* 0xe51a */
            {8'h00}, /* 0xe519 */
            {8'h00}, /* 0xe518 */
            {8'h00}, /* 0xe517 */
            {8'h00}, /* 0xe516 */
            {8'h00}, /* 0xe515 */
            {8'h00}, /* 0xe514 */
            {8'h00}, /* 0xe513 */
            {8'h00}, /* 0xe512 */
            {8'h00}, /* 0xe511 */
            {8'h00}, /* 0xe510 */
            {8'h00}, /* 0xe50f */
            {8'h00}, /* 0xe50e */
            {8'h00}, /* 0xe50d */
            {8'h00}, /* 0xe50c */
            {8'h00}, /* 0xe50b */
            {8'h00}, /* 0xe50a */
            {8'h00}, /* 0xe509 */
            {8'h00}, /* 0xe508 */
            {8'h00}, /* 0xe507 */
            {8'h00}, /* 0xe506 */
            {8'h00}, /* 0xe505 */
            {8'h00}, /* 0xe504 */
            {8'h00}, /* 0xe503 */
            {8'h00}, /* 0xe502 */
            {8'h00}, /* 0xe501 */
            {8'h00}, /* 0xe500 */
            {8'h00}, /* 0xe4ff */
            {8'h00}, /* 0xe4fe */
            {8'h00}, /* 0xe4fd */
            {8'h00}, /* 0xe4fc */
            {8'h00}, /* 0xe4fb */
            {8'h00}, /* 0xe4fa */
            {8'h00}, /* 0xe4f9 */
            {8'h00}, /* 0xe4f8 */
            {8'h00}, /* 0xe4f7 */
            {8'h00}, /* 0xe4f6 */
            {8'h00}, /* 0xe4f5 */
            {8'h00}, /* 0xe4f4 */
            {8'h00}, /* 0xe4f3 */
            {8'h00}, /* 0xe4f2 */
            {8'h00}, /* 0xe4f1 */
            {8'h00}, /* 0xe4f0 */
            {8'h00}, /* 0xe4ef */
            {8'h00}, /* 0xe4ee */
            {8'h00}, /* 0xe4ed */
            {8'h00}, /* 0xe4ec */
            {8'h00}, /* 0xe4eb */
            {8'h00}, /* 0xe4ea */
            {8'h00}, /* 0xe4e9 */
            {8'h00}, /* 0xe4e8 */
            {8'h00}, /* 0xe4e7 */
            {8'h00}, /* 0xe4e6 */
            {8'h00}, /* 0xe4e5 */
            {8'h00}, /* 0xe4e4 */
            {8'h00}, /* 0xe4e3 */
            {8'h00}, /* 0xe4e2 */
            {8'h00}, /* 0xe4e1 */
            {8'h00}, /* 0xe4e0 */
            {8'h00}, /* 0xe4df */
            {8'h00}, /* 0xe4de */
            {8'h00}, /* 0xe4dd */
            {8'h00}, /* 0xe4dc */
            {8'h00}, /* 0xe4db */
            {8'h00}, /* 0xe4da */
            {8'h00}, /* 0xe4d9 */
            {8'h00}, /* 0xe4d8 */
            {8'h00}, /* 0xe4d7 */
            {8'h00}, /* 0xe4d6 */
            {8'h00}, /* 0xe4d5 */
            {8'h00}, /* 0xe4d4 */
            {8'h00}, /* 0xe4d3 */
            {8'h00}, /* 0xe4d2 */
            {8'h00}, /* 0xe4d1 */
            {8'h00}, /* 0xe4d0 */
            {8'h00}, /* 0xe4cf */
            {8'h00}, /* 0xe4ce */
            {8'h00}, /* 0xe4cd */
            {8'h00}, /* 0xe4cc */
            {8'h00}, /* 0xe4cb */
            {8'h00}, /* 0xe4ca */
            {8'h00}, /* 0xe4c9 */
            {8'h00}, /* 0xe4c8 */
            {8'h00}, /* 0xe4c7 */
            {8'h00}, /* 0xe4c6 */
            {8'h00}, /* 0xe4c5 */
            {8'h00}, /* 0xe4c4 */
            {8'h00}, /* 0xe4c3 */
            {8'h00}, /* 0xe4c2 */
            {8'h00}, /* 0xe4c1 */
            {8'h00}, /* 0xe4c0 */
            {8'h00}, /* 0xe4bf */
            {8'h00}, /* 0xe4be */
            {8'h00}, /* 0xe4bd */
            {8'h00}, /* 0xe4bc */
            {8'h00}, /* 0xe4bb */
            {8'h00}, /* 0xe4ba */
            {8'h00}, /* 0xe4b9 */
            {8'h00}, /* 0xe4b8 */
            {8'h00}, /* 0xe4b7 */
            {8'h00}, /* 0xe4b6 */
            {8'h00}, /* 0xe4b5 */
            {8'h00}, /* 0xe4b4 */
            {8'h00}, /* 0xe4b3 */
            {8'h00}, /* 0xe4b2 */
            {8'h00}, /* 0xe4b1 */
            {8'h00}, /* 0xe4b0 */
            {8'h00}, /* 0xe4af */
            {8'h00}, /* 0xe4ae */
            {8'h00}, /* 0xe4ad */
            {8'h00}, /* 0xe4ac */
            {8'h00}, /* 0xe4ab */
            {8'h00}, /* 0xe4aa */
            {8'h00}, /* 0xe4a9 */
            {8'h00}, /* 0xe4a8 */
            {8'h00}, /* 0xe4a7 */
            {8'h00}, /* 0xe4a6 */
            {8'h00}, /* 0xe4a5 */
            {8'h00}, /* 0xe4a4 */
            {8'h00}, /* 0xe4a3 */
            {8'h00}, /* 0xe4a2 */
            {8'h00}, /* 0xe4a1 */
            {8'h00}, /* 0xe4a0 */
            {8'h00}, /* 0xe49f */
            {8'h00}, /* 0xe49e */
            {8'h00}, /* 0xe49d */
            {8'h00}, /* 0xe49c */
            {8'h00}, /* 0xe49b */
            {8'h00}, /* 0xe49a */
            {8'h00}, /* 0xe499 */
            {8'h00}, /* 0xe498 */
            {8'h00}, /* 0xe497 */
            {8'h00}, /* 0xe496 */
            {8'h00}, /* 0xe495 */
            {8'h00}, /* 0xe494 */
            {8'h00}, /* 0xe493 */
            {8'h00}, /* 0xe492 */
            {8'h00}, /* 0xe491 */
            {8'h00}, /* 0xe490 */
            {8'h00}, /* 0xe48f */
            {8'h00}, /* 0xe48e */
            {8'h00}, /* 0xe48d */
            {8'h00}, /* 0xe48c */
            {8'h00}, /* 0xe48b */
            {8'h00}, /* 0xe48a */
            {8'h00}, /* 0xe489 */
            {8'h00}, /* 0xe488 */
            {8'h00}, /* 0xe487 */
            {8'h00}, /* 0xe486 */
            {8'h00}, /* 0xe485 */
            {8'h00}, /* 0xe484 */
            {8'h00}, /* 0xe483 */
            {8'h00}, /* 0xe482 */
            {8'h00}, /* 0xe481 */
            {8'h00}, /* 0xe480 */
            {8'h00}, /* 0xe47f */
            {8'h00}, /* 0xe47e */
            {8'h00}, /* 0xe47d */
            {8'h00}, /* 0xe47c */
            {8'h00}, /* 0xe47b */
            {8'h00}, /* 0xe47a */
            {8'h00}, /* 0xe479 */
            {8'h00}, /* 0xe478 */
            {8'h00}, /* 0xe477 */
            {8'h00}, /* 0xe476 */
            {8'h00}, /* 0xe475 */
            {8'h00}, /* 0xe474 */
            {8'h00}, /* 0xe473 */
            {8'h00}, /* 0xe472 */
            {8'h00}, /* 0xe471 */
            {8'h00}, /* 0xe470 */
            {8'h00}, /* 0xe46f */
            {8'h00}, /* 0xe46e */
            {8'h00}, /* 0xe46d */
            {8'h00}, /* 0xe46c */
            {8'h00}, /* 0xe46b */
            {8'h00}, /* 0xe46a */
            {8'h00}, /* 0xe469 */
            {8'h00}, /* 0xe468 */
            {8'h00}, /* 0xe467 */
            {8'h00}, /* 0xe466 */
            {8'h00}, /* 0xe465 */
            {8'h00}, /* 0xe464 */
            {8'h00}, /* 0xe463 */
            {8'h00}, /* 0xe462 */
            {8'h00}, /* 0xe461 */
            {8'h00}, /* 0xe460 */
            {8'h00}, /* 0xe45f */
            {8'h00}, /* 0xe45e */
            {8'h00}, /* 0xe45d */
            {8'h00}, /* 0xe45c */
            {8'h00}, /* 0xe45b */
            {8'h00}, /* 0xe45a */
            {8'h00}, /* 0xe459 */
            {8'h00}, /* 0xe458 */
            {8'h00}, /* 0xe457 */
            {8'h00}, /* 0xe456 */
            {8'h00}, /* 0xe455 */
            {8'h00}, /* 0xe454 */
            {8'h00}, /* 0xe453 */
            {8'h00}, /* 0xe452 */
            {8'h00}, /* 0xe451 */
            {8'h00}, /* 0xe450 */
            {8'h00}, /* 0xe44f */
            {8'h00}, /* 0xe44e */
            {8'h00}, /* 0xe44d */
            {8'h00}, /* 0xe44c */
            {8'h00}, /* 0xe44b */
            {8'h00}, /* 0xe44a */
            {8'h00}, /* 0xe449 */
            {8'h00}, /* 0xe448 */
            {8'h00}, /* 0xe447 */
            {8'h00}, /* 0xe446 */
            {8'h00}, /* 0xe445 */
            {8'h00}, /* 0xe444 */
            {8'h00}, /* 0xe443 */
            {8'h00}, /* 0xe442 */
            {8'h00}, /* 0xe441 */
            {8'h00}, /* 0xe440 */
            {8'h00}, /* 0xe43f */
            {8'h00}, /* 0xe43e */
            {8'h00}, /* 0xe43d */
            {8'h00}, /* 0xe43c */
            {8'h00}, /* 0xe43b */
            {8'h00}, /* 0xe43a */
            {8'h00}, /* 0xe439 */
            {8'h00}, /* 0xe438 */
            {8'h00}, /* 0xe437 */
            {8'h00}, /* 0xe436 */
            {8'h00}, /* 0xe435 */
            {8'h00}, /* 0xe434 */
            {8'h00}, /* 0xe433 */
            {8'h00}, /* 0xe432 */
            {8'h00}, /* 0xe431 */
            {8'h00}, /* 0xe430 */
            {8'h00}, /* 0xe42f */
            {8'h00}, /* 0xe42e */
            {8'h00}, /* 0xe42d */
            {8'h00}, /* 0xe42c */
            {8'h00}, /* 0xe42b */
            {8'h00}, /* 0xe42a */
            {8'h00}, /* 0xe429 */
            {8'h00}, /* 0xe428 */
            {8'h00}, /* 0xe427 */
            {8'h00}, /* 0xe426 */
            {8'h00}, /* 0xe425 */
            {8'h00}, /* 0xe424 */
            {8'h00}, /* 0xe423 */
            {8'h00}, /* 0xe422 */
            {8'h00}, /* 0xe421 */
            {8'h00}, /* 0xe420 */
            {8'h00}, /* 0xe41f */
            {8'h00}, /* 0xe41e */
            {8'h00}, /* 0xe41d */
            {8'h00}, /* 0xe41c */
            {8'h00}, /* 0xe41b */
            {8'h00}, /* 0xe41a */
            {8'h00}, /* 0xe419 */
            {8'h00}, /* 0xe418 */
            {8'h00}, /* 0xe417 */
            {8'h00}, /* 0xe416 */
            {8'h00}, /* 0xe415 */
            {8'h00}, /* 0xe414 */
            {8'h00}, /* 0xe413 */
            {8'h00}, /* 0xe412 */
            {8'h00}, /* 0xe411 */
            {8'h00}, /* 0xe410 */
            {8'h00}, /* 0xe40f */
            {8'h00}, /* 0xe40e */
            {8'h00}, /* 0xe40d */
            {8'h00}, /* 0xe40c */
            {8'h00}, /* 0xe40b */
            {8'h00}, /* 0xe40a */
            {8'h00}, /* 0xe409 */
            {8'h00}, /* 0xe408 */
            {8'h00}, /* 0xe407 */
            {8'h00}, /* 0xe406 */
            {8'h00}, /* 0xe405 */
            {8'h00}, /* 0xe404 */
            {8'h00}, /* 0xe403 */
            {8'h00}, /* 0xe402 */
            {8'h00}, /* 0xe401 */
            {8'h00}, /* 0xe400 */
            {8'h00}, /* 0xe3ff */
            {8'h00}, /* 0xe3fe */
            {8'h00}, /* 0xe3fd */
            {8'h00}, /* 0xe3fc */
            {8'h00}, /* 0xe3fb */
            {8'h00}, /* 0xe3fa */
            {8'h00}, /* 0xe3f9 */
            {8'h00}, /* 0xe3f8 */
            {8'h00}, /* 0xe3f7 */
            {8'h00}, /* 0xe3f6 */
            {8'h00}, /* 0xe3f5 */
            {8'h00}, /* 0xe3f4 */
            {8'h00}, /* 0xe3f3 */
            {8'h00}, /* 0xe3f2 */
            {8'h00}, /* 0xe3f1 */
            {8'h00}, /* 0xe3f0 */
            {8'h00}, /* 0xe3ef */
            {8'h00}, /* 0xe3ee */
            {8'h00}, /* 0xe3ed */
            {8'h00}, /* 0xe3ec */
            {8'h00}, /* 0xe3eb */
            {8'h00}, /* 0xe3ea */
            {8'h00}, /* 0xe3e9 */
            {8'h00}, /* 0xe3e8 */
            {8'h00}, /* 0xe3e7 */
            {8'h00}, /* 0xe3e6 */
            {8'h00}, /* 0xe3e5 */
            {8'h00}, /* 0xe3e4 */
            {8'h00}, /* 0xe3e3 */
            {8'h00}, /* 0xe3e2 */
            {8'h00}, /* 0xe3e1 */
            {8'h00}, /* 0xe3e0 */
            {8'h00}, /* 0xe3df */
            {8'h00}, /* 0xe3de */
            {8'h00}, /* 0xe3dd */
            {8'h00}, /* 0xe3dc */
            {8'h00}, /* 0xe3db */
            {8'h00}, /* 0xe3da */
            {8'h00}, /* 0xe3d9 */
            {8'h00}, /* 0xe3d8 */
            {8'h00}, /* 0xe3d7 */
            {8'h00}, /* 0xe3d6 */
            {8'h00}, /* 0xe3d5 */
            {8'h00}, /* 0xe3d4 */
            {8'h00}, /* 0xe3d3 */
            {8'h00}, /* 0xe3d2 */
            {8'h00}, /* 0xe3d1 */
            {8'h00}, /* 0xe3d0 */
            {8'h00}, /* 0xe3cf */
            {8'h00}, /* 0xe3ce */
            {8'h00}, /* 0xe3cd */
            {8'h00}, /* 0xe3cc */
            {8'h00}, /* 0xe3cb */
            {8'h00}, /* 0xe3ca */
            {8'h00}, /* 0xe3c9 */
            {8'h00}, /* 0xe3c8 */
            {8'h00}, /* 0xe3c7 */
            {8'h00}, /* 0xe3c6 */
            {8'h00}, /* 0xe3c5 */
            {8'h00}, /* 0xe3c4 */
            {8'h00}, /* 0xe3c3 */
            {8'h00}, /* 0xe3c2 */
            {8'h00}, /* 0xe3c1 */
            {8'h00}, /* 0xe3c0 */
            {8'h00}, /* 0xe3bf */
            {8'h00}, /* 0xe3be */
            {8'h00}, /* 0xe3bd */
            {8'h00}, /* 0xe3bc */
            {8'h00}, /* 0xe3bb */
            {8'h00}, /* 0xe3ba */
            {8'h00}, /* 0xe3b9 */
            {8'h00}, /* 0xe3b8 */
            {8'h00}, /* 0xe3b7 */
            {8'h00}, /* 0xe3b6 */
            {8'h00}, /* 0xe3b5 */
            {8'h00}, /* 0xe3b4 */
            {8'h00}, /* 0xe3b3 */
            {8'h00}, /* 0xe3b2 */
            {8'h00}, /* 0xe3b1 */
            {8'h00}, /* 0xe3b0 */
            {8'h00}, /* 0xe3af */
            {8'h00}, /* 0xe3ae */
            {8'h00}, /* 0xe3ad */
            {8'h00}, /* 0xe3ac */
            {8'h00}, /* 0xe3ab */
            {8'h00}, /* 0xe3aa */
            {8'h00}, /* 0xe3a9 */
            {8'h00}, /* 0xe3a8 */
            {8'h00}, /* 0xe3a7 */
            {8'h00}, /* 0xe3a6 */
            {8'h00}, /* 0xe3a5 */
            {8'h00}, /* 0xe3a4 */
            {8'h00}, /* 0xe3a3 */
            {8'h00}, /* 0xe3a2 */
            {8'h00}, /* 0xe3a1 */
            {8'h00}, /* 0xe3a0 */
            {8'h00}, /* 0xe39f */
            {8'h00}, /* 0xe39e */
            {8'h00}, /* 0xe39d */
            {8'h00}, /* 0xe39c */
            {8'h00}, /* 0xe39b */
            {8'h00}, /* 0xe39a */
            {8'h00}, /* 0xe399 */
            {8'h00}, /* 0xe398 */
            {8'h00}, /* 0xe397 */
            {8'h00}, /* 0xe396 */
            {8'h00}, /* 0xe395 */
            {8'h00}, /* 0xe394 */
            {8'h00}, /* 0xe393 */
            {8'h00}, /* 0xe392 */
            {8'h00}, /* 0xe391 */
            {8'h00}, /* 0xe390 */
            {8'h00}, /* 0xe38f */
            {8'h00}, /* 0xe38e */
            {8'h00}, /* 0xe38d */
            {8'h00}, /* 0xe38c */
            {8'h00}, /* 0xe38b */
            {8'h00}, /* 0xe38a */
            {8'h00}, /* 0xe389 */
            {8'h00}, /* 0xe388 */
            {8'h00}, /* 0xe387 */
            {8'h00}, /* 0xe386 */
            {8'h00}, /* 0xe385 */
            {8'h00}, /* 0xe384 */
            {8'h00}, /* 0xe383 */
            {8'h00}, /* 0xe382 */
            {8'h00}, /* 0xe381 */
            {8'h00}, /* 0xe380 */
            {8'h00}, /* 0xe37f */
            {8'h00}, /* 0xe37e */
            {8'h00}, /* 0xe37d */
            {8'h00}, /* 0xe37c */
            {8'h00}, /* 0xe37b */
            {8'h00}, /* 0xe37a */
            {8'h00}, /* 0xe379 */
            {8'h00}, /* 0xe378 */
            {8'h00}, /* 0xe377 */
            {8'h00}, /* 0xe376 */
            {8'h00}, /* 0xe375 */
            {8'h00}, /* 0xe374 */
            {8'h00}, /* 0xe373 */
            {8'h00}, /* 0xe372 */
            {8'h00}, /* 0xe371 */
            {8'h00}, /* 0xe370 */
            {8'h00}, /* 0xe36f */
            {8'h00}, /* 0xe36e */
            {8'h00}, /* 0xe36d */
            {8'h00}, /* 0xe36c */
            {8'h00}, /* 0xe36b */
            {8'h00}, /* 0xe36a */
            {8'h00}, /* 0xe369 */
            {8'h00}, /* 0xe368 */
            {8'h00}, /* 0xe367 */
            {8'h00}, /* 0xe366 */
            {8'h00}, /* 0xe365 */
            {8'h00}, /* 0xe364 */
            {8'h00}, /* 0xe363 */
            {8'h00}, /* 0xe362 */
            {8'h00}, /* 0xe361 */
            {8'h00}, /* 0xe360 */
            {8'h00}, /* 0xe35f */
            {8'h00}, /* 0xe35e */
            {8'h00}, /* 0xe35d */
            {8'h00}, /* 0xe35c */
            {8'h00}, /* 0xe35b */
            {8'h00}, /* 0xe35a */
            {8'h00}, /* 0xe359 */
            {8'h00}, /* 0xe358 */
            {8'h00}, /* 0xe357 */
            {8'h00}, /* 0xe356 */
            {8'h00}, /* 0xe355 */
            {8'h00}, /* 0xe354 */
            {8'h00}, /* 0xe353 */
            {8'h00}, /* 0xe352 */
            {8'h00}, /* 0xe351 */
            {8'h00}, /* 0xe350 */
            {8'h00}, /* 0xe34f */
            {8'h00}, /* 0xe34e */
            {8'h00}, /* 0xe34d */
            {8'h00}, /* 0xe34c */
            {8'h00}, /* 0xe34b */
            {8'h00}, /* 0xe34a */
            {8'h00}, /* 0xe349 */
            {8'h00}, /* 0xe348 */
            {8'h00}, /* 0xe347 */
            {8'h00}, /* 0xe346 */
            {8'h00}, /* 0xe345 */
            {8'h00}, /* 0xe344 */
            {8'h00}, /* 0xe343 */
            {8'h00}, /* 0xe342 */
            {8'h00}, /* 0xe341 */
            {8'h00}, /* 0xe340 */
            {8'h00}, /* 0xe33f */
            {8'h00}, /* 0xe33e */
            {8'h00}, /* 0xe33d */
            {8'h00}, /* 0xe33c */
            {8'h00}, /* 0xe33b */
            {8'h00}, /* 0xe33a */
            {8'h00}, /* 0xe339 */
            {8'h00}, /* 0xe338 */
            {8'h00}, /* 0xe337 */
            {8'h00}, /* 0xe336 */
            {8'h00}, /* 0xe335 */
            {8'h00}, /* 0xe334 */
            {8'h00}, /* 0xe333 */
            {8'h00}, /* 0xe332 */
            {8'h00}, /* 0xe331 */
            {8'h00}, /* 0xe330 */
            {8'h00}, /* 0xe32f */
            {8'h00}, /* 0xe32e */
            {8'h00}, /* 0xe32d */
            {8'h00}, /* 0xe32c */
            {8'h00}, /* 0xe32b */
            {8'h00}, /* 0xe32a */
            {8'h00}, /* 0xe329 */
            {8'h00}, /* 0xe328 */
            {8'h00}, /* 0xe327 */
            {8'h00}, /* 0xe326 */
            {8'h00}, /* 0xe325 */
            {8'h00}, /* 0xe324 */
            {8'h00}, /* 0xe323 */
            {8'h00}, /* 0xe322 */
            {8'h00}, /* 0xe321 */
            {8'h00}, /* 0xe320 */
            {8'h00}, /* 0xe31f */
            {8'h00}, /* 0xe31e */
            {8'h00}, /* 0xe31d */
            {8'h00}, /* 0xe31c */
            {8'h00}, /* 0xe31b */
            {8'h00}, /* 0xe31a */
            {8'h00}, /* 0xe319 */
            {8'h00}, /* 0xe318 */
            {8'h00}, /* 0xe317 */
            {8'h00}, /* 0xe316 */
            {8'h00}, /* 0xe315 */
            {8'h00}, /* 0xe314 */
            {8'h00}, /* 0xe313 */
            {8'h00}, /* 0xe312 */
            {8'h00}, /* 0xe311 */
            {8'h00}, /* 0xe310 */
            {8'h00}, /* 0xe30f */
            {8'h00}, /* 0xe30e */
            {8'h00}, /* 0xe30d */
            {8'h00}, /* 0xe30c */
            {8'h00}, /* 0xe30b */
            {8'h00}, /* 0xe30a */
            {8'h00}, /* 0xe309 */
            {8'h00}, /* 0xe308 */
            {8'h00}, /* 0xe307 */
            {8'h00}, /* 0xe306 */
            {8'h00}, /* 0xe305 */
            {8'h00}, /* 0xe304 */
            {8'h00}, /* 0xe303 */
            {8'h00}, /* 0xe302 */
            {8'h00}, /* 0xe301 */
            {8'h00}, /* 0xe300 */
            {8'h00}, /* 0xe2ff */
            {8'h00}, /* 0xe2fe */
            {8'h00}, /* 0xe2fd */
            {8'h00}, /* 0xe2fc */
            {8'h00}, /* 0xe2fb */
            {8'h00}, /* 0xe2fa */
            {8'h00}, /* 0xe2f9 */
            {8'h00}, /* 0xe2f8 */
            {8'h00}, /* 0xe2f7 */
            {8'h00}, /* 0xe2f6 */
            {8'h00}, /* 0xe2f5 */
            {8'h00}, /* 0xe2f4 */
            {8'h00}, /* 0xe2f3 */
            {8'h00}, /* 0xe2f2 */
            {8'h00}, /* 0xe2f1 */
            {8'h00}, /* 0xe2f0 */
            {8'h00}, /* 0xe2ef */
            {8'h00}, /* 0xe2ee */
            {8'h00}, /* 0xe2ed */
            {8'h00}, /* 0xe2ec */
            {8'h00}, /* 0xe2eb */
            {8'h00}, /* 0xe2ea */
            {8'h00}, /* 0xe2e9 */
            {8'h00}, /* 0xe2e8 */
            {8'h00}, /* 0xe2e7 */
            {8'h00}, /* 0xe2e6 */
            {8'h00}, /* 0xe2e5 */
            {8'h00}, /* 0xe2e4 */
            {8'h00}, /* 0xe2e3 */
            {8'h00}, /* 0xe2e2 */
            {8'h00}, /* 0xe2e1 */
            {8'h00}, /* 0xe2e0 */
            {8'h00}, /* 0xe2df */
            {8'h00}, /* 0xe2de */
            {8'h00}, /* 0xe2dd */
            {8'h00}, /* 0xe2dc */
            {8'h00}, /* 0xe2db */
            {8'h00}, /* 0xe2da */
            {8'h00}, /* 0xe2d9 */
            {8'h00}, /* 0xe2d8 */
            {8'h00}, /* 0xe2d7 */
            {8'h00}, /* 0xe2d6 */
            {8'h00}, /* 0xe2d5 */
            {8'h00}, /* 0xe2d4 */
            {8'h00}, /* 0xe2d3 */
            {8'h00}, /* 0xe2d2 */
            {8'h00}, /* 0xe2d1 */
            {8'h00}, /* 0xe2d0 */
            {8'h00}, /* 0xe2cf */
            {8'h00}, /* 0xe2ce */
            {8'h00}, /* 0xe2cd */
            {8'h00}, /* 0xe2cc */
            {8'h00}, /* 0xe2cb */
            {8'h00}, /* 0xe2ca */
            {8'h00}, /* 0xe2c9 */
            {8'h00}, /* 0xe2c8 */
            {8'h00}, /* 0xe2c7 */
            {8'h00}, /* 0xe2c6 */
            {8'h00}, /* 0xe2c5 */
            {8'h00}, /* 0xe2c4 */
            {8'h00}, /* 0xe2c3 */
            {8'h00}, /* 0xe2c2 */
            {8'h00}, /* 0xe2c1 */
            {8'h00}, /* 0xe2c0 */
            {8'h00}, /* 0xe2bf */
            {8'h00}, /* 0xe2be */
            {8'h00}, /* 0xe2bd */
            {8'h00}, /* 0xe2bc */
            {8'h00}, /* 0xe2bb */
            {8'h00}, /* 0xe2ba */
            {8'h00}, /* 0xe2b9 */
            {8'h00}, /* 0xe2b8 */
            {8'h00}, /* 0xe2b7 */
            {8'h00}, /* 0xe2b6 */
            {8'h00}, /* 0xe2b5 */
            {8'h00}, /* 0xe2b4 */
            {8'h00}, /* 0xe2b3 */
            {8'h00}, /* 0xe2b2 */
            {8'h00}, /* 0xe2b1 */
            {8'h00}, /* 0xe2b0 */
            {8'h00}, /* 0xe2af */
            {8'h00}, /* 0xe2ae */
            {8'h00}, /* 0xe2ad */
            {8'h00}, /* 0xe2ac */
            {8'h00}, /* 0xe2ab */
            {8'h00}, /* 0xe2aa */
            {8'h00}, /* 0xe2a9 */
            {8'h00}, /* 0xe2a8 */
            {8'h00}, /* 0xe2a7 */
            {8'h00}, /* 0xe2a6 */
            {8'h00}, /* 0xe2a5 */
            {8'h00}, /* 0xe2a4 */
            {8'h00}, /* 0xe2a3 */
            {8'h00}, /* 0xe2a2 */
            {8'h00}, /* 0xe2a1 */
            {8'h00}, /* 0xe2a0 */
            {8'h00}, /* 0xe29f */
            {8'h00}, /* 0xe29e */
            {8'h00}, /* 0xe29d */
            {8'h00}, /* 0xe29c */
            {8'h00}, /* 0xe29b */
            {8'h00}, /* 0xe29a */
            {8'h00}, /* 0xe299 */
            {8'h00}, /* 0xe298 */
            {8'h00}, /* 0xe297 */
            {8'h00}, /* 0xe296 */
            {8'h00}, /* 0xe295 */
            {8'h00}, /* 0xe294 */
            {8'h00}, /* 0xe293 */
            {8'h00}, /* 0xe292 */
            {8'h00}, /* 0xe291 */
            {8'h00}, /* 0xe290 */
            {8'h00}, /* 0xe28f */
            {8'h00}, /* 0xe28e */
            {8'h00}, /* 0xe28d */
            {8'h00}, /* 0xe28c */
            {8'h00}, /* 0xe28b */
            {8'h00}, /* 0xe28a */
            {8'h00}, /* 0xe289 */
            {8'h00}, /* 0xe288 */
            {8'h00}, /* 0xe287 */
            {8'h00}, /* 0xe286 */
            {8'h00}, /* 0xe285 */
            {8'h00}, /* 0xe284 */
            {8'h00}, /* 0xe283 */
            {8'h00}, /* 0xe282 */
            {8'h00}, /* 0xe281 */
            {8'h00}, /* 0xe280 */
            {8'h00}, /* 0xe27f */
            {8'h00}, /* 0xe27e */
            {8'h00}, /* 0xe27d */
            {8'h00}, /* 0xe27c */
            {8'h00}, /* 0xe27b */
            {8'h00}, /* 0xe27a */
            {8'h00}, /* 0xe279 */
            {8'h00}, /* 0xe278 */
            {8'h00}, /* 0xe277 */
            {8'h00}, /* 0xe276 */
            {8'h00}, /* 0xe275 */
            {8'h00}, /* 0xe274 */
            {8'h00}, /* 0xe273 */
            {8'h00}, /* 0xe272 */
            {8'h00}, /* 0xe271 */
            {8'h00}, /* 0xe270 */
            {8'h00}, /* 0xe26f */
            {8'h00}, /* 0xe26e */
            {8'h00}, /* 0xe26d */
            {8'h00}, /* 0xe26c */
            {8'h00}, /* 0xe26b */
            {8'h00}, /* 0xe26a */
            {8'h00}, /* 0xe269 */
            {8'h00}, /* 0xe268 */
            {8'h00}, /* 0xe267 */
            {8'h00}, /* 0xe266 */
            {8'h00}, /* 0xe265 */
            {8'h00}, /* 0xe264 */
            {8'h00}, /* 0xe263 */
            {8'h00}, /* 0xe262 */
            {8'h00}, /* 0xe261 */
            {8'h00}, /* 0xe260 */
            {8'h00}, /* 0xe25f */
            {8'h00}, /* 0xe25e */
            {8'h00}, /* 0xe25d */
            {8'h00}, /* 0xe25c */
            {8'h00}, /* 0xe25b */
            {8'h00}, /* 0xe25a */
            {8'h00}, /* 0xe259 */
            {8'h00}, /* 0xe258 */
            {8'h00}, /* 0xe257 */
            {8'h00}, /* 0xe256 */
            {8'h00}, /* 0xe255 */
            {8'h00}, /* 0xe254 */
            {8'h00}, /* 0xe253 */
            {8'h00}, /* 0xe252 */
            {8'h00}, /* 0xe251 */
            {8'h00}, /* 0xe250 */
            {8'h00}, /* 0xe24f */
            {8'h00}, /* 0xe24e */
            {8'h00}, /* 0xe24d */
            {8'h00}, /* 0xe24c */
            {8'h00}, /* 0xe24b */
            {8'h00}, /* 0xe24a */
            {8'h00}, /* 0xe249 */
            {8'h00}, /* 0xe248 */
            {8'h00}, /* 0xe247 */
            {8'h00}, /* 0xe246 */
            {8'h00}, /* 0xe245 */
            {8'h00}, /* 0xe244 */
            {8'h00}, /* 0xe243 */
            {8'h00}, /* 0xe242 */
            {8'h00}, /* 0xe241 */
            {8'h00}, /* 0xe240 */
            {8'h00}, /* 0xe23f */
            {8'h00}, /* 0xe23e */
            {8'h00}, /* 0xe23d */
            {8'h00}, /* 0xe23c */
            {8'h00}, /* 0xe23b */
            {8'h00}, /* 0xe23a */
            {8'h00}, /* 0xe239 */
            {8'h00}, /* 0xe238 */
            {8'h00}, /* 0xe237 */
            {8'h00}, /* 0xe236 */
            {8'h00}, /* 0xe235 */
            {8'h00}, /* 0xe234 */
            {8'h00}, /* 0xe233 */
            {8'h00}, /* 0xe232 */
            {8'h00}, /* 0xe231 */
            {8'h00}, /* 0xe230 */
            {8'h00}, /* 0xe22f */
            {8'h00}, /* 0xe22e */
            {8'h00}, /* 0xe22d */
            {8'h00}, /* 0xe22c */
            {8'h00}, /* 0xe22b */
            {8'h00}, /* 0xe22a */
            {8'h00}, /* 0xe229 */
            {8'h00}, /* 0xe228 */
            {8'h00}, /* 0xe227 */
            {8'h00}, /* 0xe226 */
            {8'h00}, /* 0xe225 */
            {8'h00}, /* 0xe224 */
            {8'h00}, /* 0xe223 */
            {8'h00}, /* 0xe222 */
            {8'h00}, /* 0xe221 */
            {8'h00}, /* 0xe220 */
            {8'h00}, /* 0xe21f */
            {8'h00}, /* 0xe21e */
            {8'h00}, /* 0xe21d */
            {8'h00}, /* 0xe21c */
            {8'h00}, /* 0xe21b */
            {8'h00}, /* 0xe21a */
            {8'h00}, /* 0xe219 */
            {8'h00}, /* 0xe218 */
            {8'h00}, /* 0xe217 */
            {8'h00}, /* 0xe216 */
            {8'h00}, /* 0xe215 */
            {8'h00}, /* 0xe214 */
            {8'h00}, /* 0xe213 */
            {8'h00}, /* 0xe212 */
            {8'h00}, /* 0xe211 */
            {8'h00}, /* 0xe210 */
            {8'h00}, /* 0xe20f */
            {8'h00}, /* 0xe20e */
            {8'h00}, /* 0xe20d */
            {8'h00}, /* 0xe20c */
            {8'h00}, /* 0xe20b */
            {8'h00}, /* 0xe20a */
            {8'h00}, /* 0xe209 */
            {8'h00}, /* 0xe208 */
            {8'h00}, /* 0xe207 */
            {8'h00}, /* 0xe206 */
            {8'h00}, /* 0xe205 */
            {8'h00}, /* 0xe204 */
            {8'h00}, /* 0xe203 */
            {8'h00}, /* 0xe202 */
            {8'h00}, /* 0xe201 */
            {8'h00}, /* 0xe200 */
            {8'h00}, /* 0xe1ff */
            {8'h00}, /* 0xe1fe */
            {8'h00}, /* 0xe1fd */
            {8'h00}, /* 0xe1fc */
            {8'h00}, /* 0xe1fb */
            {8'h00}, /* 0xe1fa */
            {8'h00}, /* 0xe1f9 */
            {8'h00}, /* 0xe1f8 */
            {8'h00}, /* 0xe1f7 */
            {8'h00}, /* 0xe1f6 */
            {8'h00}, /* 0xe1f5 */
            {8'h00}, /* 0xe1f4 */
            {8'h00}, /* 0xe1f3 */
            {8'h00}, /* 0xe1f2 */
            {8'h00}, /* 0xe1f1 */
            {8'h00}, /* 0xe1f0 */
            {8'h00}, /* 0xe1ef */
            {8'h00}, /* 0xe1ee */
            {8'h00}, /* 0xe1ed */
            {8'h00}, /* 0xe1ec */
            {8'h00}, /* 0xe1eb */
            {8'h00}, /* 0xe1ea */
            {8'h00}, /* 0xe1e9 */
            {8'h00}, /* 0xe1e8 */
            {8'h00}, /* 0xe1e7 */
            {8'h00}, /* 0xe1e6 */
            {8'h00}, /* 0xe1e5 */
            {8'h00}, /* 0xe1e4 */
            {8'h00}, /* 0xe1e3 */
            {8'h00}, /* 0xe1e2 */
            {8'h00}, /* 0xe1e1 */
            {8'h00}, /* 0xe1e0 */
            {8'h00}, /* 0xe1df */
            {8'h00}, /* 0xe1de */
            {8'h00}, /* 0xe1dd */
            {8'h00}, /* 0xe1dc */
            {8'h00}, /* 0xe1db */
            {8'h00}, /* 0xe1da */
            {8'h00}, /* 0xe1d9 */
            {8'h00}, /* 0xe1d8 */
            {8'h00}, /* 0xe1d7 */
            {8'h00}, /* 0xe1d6 */
            {8'h00}, /* 0xe1d5 */
            {8'h00}, /* 0xe1d4 */
            {8'h00}, /* 0xe1d3 */
            {8'h00}, /* 0xe1d2 */
            {8'h00}, /* 0xe1d1 */
            {8'h00}, /* 0xe1d0 */
            {8'h00}, /* 0xe1cf */
            {8'h00}, /* 0xe1ce */
            {8'h00}, /* 0xe1cd */
            {8'h00}, /* 0xe1cc */
            {8'h00}, /* 0xe1cb */
            {8'h00}, /* 0xe1ca */
            {8'h00}, /* 0xe1c9 */
            {8'h00}, /* 0xe1c8 */
            {8'h00}, /* 0xe1c7 */
            {8'h00}, /* 0xe1c6 */
            {8'h00}, /* 0xe1c5 */
            {8'h00}, /* 0xe1c4 */
            {8'h00}, /* 0xe1c3 */
            {8'h00}, /* 0xe1c2 */
            {8'h00}, /* 0xe1c1 */
            {8'h00}, /* 0xe1c0 */
            {8'h00}, /* 0xe1bf */
            {8'h00}, /* 0xe1be */
            {8'h00}, /* 0xe1bd */
            {8'h00}, /* 0xe1bc */
            {8'h00}, /* 0xe1bb */
            {8'h00}, /* 0xe1ba */
            {8'h00}, /* 0xe1b9 */
            {8'h00}, /* 0xe1b8 */
            {8'h00}, /* 0xe1b7 */
            {8'h00}, /* 0xe1b6 */
            {8'h00}, /* 0xe1b5 */
            {8'h00}, /* 0xe1b4 */
            {8'h00}, /* 0xe1b3 */
            {8'h00}, /* 0xe1b2 */
            {8'h00}, /* 0xe1b1 */
            {8'h00}, /* 0xe1b0 */
            {8'h00}, /* 0xe1af */
            {8'h00}, /* 0xe1ae */
            {8'h00}, /* 0xe1ad */
            {8'h00}, /* 0xe1ac */
            {8'h00}, /* 0xe1ab */
            {8'h00}, /* 0xe1aa */
            {8'h00}, /* 0xe1a9 */
            {8'h00}, /* 0xe1a8 */
            {8'h00}, /* 0xe1a7 */
            {8'h00}, /* 0xe1a6 */
            {8'h00}, /* 0xe1a5 */
            {8'h00}, /* 0xe1a4 */
            {8'h00}, /* 0xe1a3 */
            {8'h00}, /* 0xe1a2 */
            {8'h00}, /* 0xe1a1 */
            {8'h00}, /* 0xe1a0 */
            {8'h00}, /* 0xe19f */
            {8'h00}, /* 0xe19e */
            {8'h00}, /* 0xe19d */
            {8'h00}, /* 0xe19c */
            {8'h00}, /* 0xe19b */
            {8'h00}, /* 0xe19a */
            {8'h00}, /* 0xe199 */
            {8'h00}, /* 0xe198 */
            {8'h00}, /* 0xe197 */
            {8'h00}, /* 0xe196 */
            {8'h00}, /* 0xe195 */
            {8'h00}, /* 0xe194 */
            {8'h00}, /* 0xe193 */
            {8'h00}, /* 0xe192 */
            {8'h00}, /* 0xe191 */
            {8'h00}, /* 0xe190 */
            {8'h00}, /* 0xe18f */
            {8'h00}, /* 0xe18e */
            {8'h00}, /* 0xe18d */
            {8'h00}, /* 0xe18c */
            {8'h00}, /* 0xe18b */
            {8'h00}, /* 0xe18a */
            {8'h00}, /* 0xe189 */
            {8'h00}, /* 0xe188 */
            {8'h00}, /* 0xe187 */
            {8'h00}, /* 0xe186 */
            {8'h00}, /* 0xe185 */
            {8'h00}, /* 0xe184 */
            {8'h00}, /* 0xe183 */
            {8'h00}, /* 0xe182 */
            {8'h00}, /* 0xe181 */
            {8'h00}, /* 0xe180 */
            {8'h00}, /* 0xe17f */
            {8'h00}, /* 0xe17e */
            {8'h00}, /* 0xe17d */
            {8'h00}, /* 0xe17c */
            {8'h00}, /* 0xe17b */
            {8'h00}, /* 0xe17a */
            {8'h00}, /* 0xe179 */
            {8'h00}, /* 0xe178 */
            {8'h00}, /* 0xe177 */
            {8'h00}, /* 0xe176 */
            {8'h00}, /* 0xe175 */
            {8'h00}, /* 0xe174 */
            {8'h00}, /* 0xe173 */
            {8'h00}, /* 0xe172 */
            {8'h00}, /* 0xe171 */
            {8'h00}, /* 0xe170 */
            {8'h00}, /* 0xe16f */
            {8'h00}, /* 0xe16e */
            {8'h00}, /* 0xe16d */
            {8'h00}, /* 0xe16c */
            {8'h00}, /* 0xe16b */
            {8'h00}, /* 0xe16a */
            {8'h00}, /* 0xe169 */
            {8'h00}, /* 0xe168 */
            {8'h00}, /* 0xe167 */
            {8'h00}, /* 0xe166 */
            {8'h00}, /* 0xe165 */
            {8'h00}, /* 0xe164 */
            {8'h00}, /* 0xe163 */
            {8'h00}, /* 0xe162 */
            {8'h00}, /* 0xe161 */
            {8'h00}, /* 0xe160 */
            {8'h00}, /* 0xe15f */
            {8'h00}, /* 0xe15e */
            {8'h00}, /* 0xe15d */
            {8'h00}, /* 0xe15c */
            {8'h00}, /* 0xe15b */
            {8'h00}, /* 0xe15a */
            {8'h00}, /* 0xe159 */
            {8'h00}, /* 0xe158 */
            {8'h00}, /* 0xe157 */
            {8'h00}, /* 0xe156 */
            {8'h00}, /* 0xe155 */
            {8'h00}, /* 0xe154 */
            {8'h00}, /* 0xe153 */
            {8'h00}, /* 0xe152 */
            {8'h00}, /* 0xe151 */
            {8'h00}, /* 0xe150 */
            {8'h00}, /* 0xe14f */
            {8'h00}, /* 0xe14e */
            {8'h00}, /* 0xe14d */
            {8'h00}, /* 0xe14c */
            {8'h00}, /* 0xe14b */
            {8'h00}, /* 0xe14a */
            {8'h00}, /* 0xe149 */
            {8'h00}, /* 0xe148 */
            {8'h00}, /* 0xe147 */
            {8'h00}, /* 0xe146 */
            {8'h00}, /* 0xe145 */
            {8'h00}, /* 0xe144 */
            {8'h00}, /* 0xe143 */
            {8'h00}, /* 0xe142 */
            {8'h00}, /* 0xe141 */
            {8'h00}, /* 0xe140 */
            {8'h00}, /* 0xe13f */
            {8'h00}, /* 0xe13e */
            {8'h00}, /* 0xe13d */
            {8'h00}, /* 0xe13c */
            {8'h00}, /* 0xe13b */
            {8'h00}, /* 0xe13a */
            {8'h00}, /* 0xe139 */
            {8'h00}, /* 0xe138 */
            {8'h00}, /* 0xe137 */
            {8'h00}, /* 0xe136 */
            {8'h00}, /* 0xe135 */
            {8'h00}, /* 0xe134 */
            {8'h00}, /* 0xe133 */
            {8'h00}, /* 0xe132 */
            {8'h00}, /* 0xe131 */
            {8'h00}, /* 0xe130 */
            {8'h00}, /* 0xe12f */
            {8'h00}, /* 0xe12e */
            {8'h00}, /* 0xe12d */
            {8'h00}, /* 0xe12c */
            {8'h00}, /* 0xe12b */
            {8'h00}, /* 0xe12a */
            {8'h00}, /* 0xe129 */
            {8'h00}, /* 0xe128 */
            {8'h00}, /* 0xe127 */
            {8'h00}, /* 0xe126 */
            {8'h00}, /* 0xe125 */
            {8'h00}, /* 0xe124 */
            {8'h00}, /* 0xe123 */
            {8'h00}, /* 0xe122 */
            {8'h00}, /* 0xe121 */
            {8'h00}, /* 0xe120 */
            {8'h00}, /* 0xe11f */
            {8'h00}, /* 0xe11e */
            {8'h00}, /* 0xe11d */
            {8'h00}, /* 0xe11c */
            {8'h00}, /* 0xe11b */
            {8'h00}, /* 0xe11a */
            {8'h00}, /* 0xe119 */
            {8'h00}, /* 0xe118 */
            {8'h00}, /* 0xe117 */
            {8'h00}, /* 0xe116 */
            {8'h00}, /* 0xe115 */
            {8'h00}, /* 0xe114 */
            {8'h00}, /* 0xe113 */
            {8'h00}, /* 0xe112 */
            {8'h00}, /* 0xe111 */
            {8'h00}, /* 0xe110 */
            {8'h00}, /* 0xe10f */
            {8'h00}, /* 0xe10e */
            {8'h00}, /* 0xe10d */
            {8'h00}, /* 0xe10c */
            {8'h00}, /* 0xe10b */
            {8'h00}, /* 0xe10a */
            {8'h00}, /* 0xe109 */
            {8'h00}, /* 0xe108 */
            {8'h00}, /* 0xe107 */
            {8'h00}, /* 0xe106 */
            {8'h00}, /* 0xe105 */
            {8'h00}, /* 0xe104 */
            {8'h00}, /* 0xe103 */
            {8'h00}, /* 0xe102 */
            {8'h00}, /* 0xe101 */
            {8'h00}, /* 0xe100 */
            {8'h00}, /* 0xe0ff */
            {8'h00}, /* 0xe0fe */
            {8'h00}, /* 0xe0fd */
            {8'h00}, /* 0xe0fc */
            {8'h00}, /* 0xe0fb */
            {8'h00}, /* 0xe0fa */
            {8'h00}, /* 0xe0f9 */
            {8'h00}, /* 0xe0f8 */
            {8'h00}, /* 0xe0f7 */
            {8'h00}, /* 0xe0f6 */
            {8'h00}, /* 0xe0f5 */
            {8'h00}, /* 0xe0f4 */
            {8'h00}, /* 0xe0f3 */
            {8'h00}, /* 0xe0f2 */
            {8'h00}, /* 0xe0f1 */
            {8'h00}, /* 0xe0f0 */
            {8'h00}, /* 0xe0ef */
            {8'h00}, /* 0xe0ee */
            {8'h00}, /* 0xe0ed */
            {8'h00}, /* 0xe0ec */
            {8'h00}, /* 0xe0eb */
            {8'h00}, /* 0xe0ea */
            {8'h00}, /* 0xe0e9 */
            {8'h00}, /* 0xe0e8 */
            {8'h00}, /* 0xe0e7 */
            {8'h00}, /* 0xe0e6 */
            {8'h00}, /* 0xe0e5 */
            {8'h00}, /* 0xe0e4 */
            {8'h00}, /* 0xe0e3 */
            {8'h00}, /* 0xe0e2 */
            {8'h00}, /* 0xe0e1 */
            {8'h00}, /* 0xe0e0 */
            {8'h00}, /* 0xe0df */
            {8'h00}, /* 0xe0de */
            {8'h00}, /* 0xe0dd */
            {8'h00}, /* 0xe0dc */
            {8'h00}, /* 0xe0db */
            {8'h00}, /* 0xe0da */
            {8'h00}, /* 0xe0d9 */
            {8'h00}, /* 0xe0d8 */
            {8'h00}, /* 0xe0d7 */
            {8'h00}, /* 0xe0d6 */
            {8'h00}, /* 0xe0d5 */
            {8'h00}, /* 0xe0d4 */
            {8'h00}, /* 0xe0d3 */
            {8'h00}, /* 0xe0d2 */
            {8'h00}, /* 0xe0d1 */
            {8'h00}, /* 0xe0d0 */
            {8'h00}, /* 0xe0cf */
            {8'h00}, /* 0xe0ce */
            {8'h00}, /* 0xe0cd */
            {8'h00}, /* 0xe0cc */
            {8'h00}, /* 0xe0cb */
            {8'h00}, /* 0xe0ca */
            {8'h00}, /* 0xe0c9 */
            {8'h00}, /* 0xe0c8 */
            {8'h00}, /* 0xe0c7 */
            {8'h00}, /* 0xe0c6 */
            {8'h00}, /* 0xe0c5 */
            {8'h00}, /* 0xe0c4 */
            {8'h00}, /* 0xe0c3 */
            {8'h00}, /* 0xe0c2 */
            {8'h00}, /* 0xe0c1 */
            {8'h00}, /* 0xe0c0 */
            {8'h00}, /* 0xe0bf */
            {8'h00}, /* 0xe0be */
            {8'h00}, /* 0xe0bd */
            {8'h00}, /* 0xe0bc */
            {8'h00}, /* 0xe0bb */
            {8'h00}, /* 0xe0ba */
            {8'h00}, /* 0xe0b9 */
            {8'h00}, /* 0xe0b8 */
            {8'h00}, /* 0xe0b7 */
            {8'h00}, /* 0xe0b6 */
            {8'h00}, /* 0xe0b5 */
            {8'h00}, /* 0xe0b4 */
            {8'h00}, /* 0xe0b3 */
            {8'h00}, /* 0xe0b2 */
            {8'h00}, /* 0xe0b1 */
            {8'h00}, /* 0xe0b0 */
            {8'h00}, /* 0xe0af */
            {8'h00}, /* 0xe0ae */
            {8'h00}, /* 0xe0ad */
            {8'h00}, /* 0xe0ac */
            {8'h00}, /* 0xe0ab */
            {8'h00}, /* 0xe0aa */
            {8'h00}, /* 0xe0a9 */
            {8'h00}, /* 0xe0a8 */
            {8'h00}, /* 0xe0a7 */
            {8'h00}, /* 0xe0a6 */
            {8'h00}, /* 0xe0a5 */
            {8'h00}, /* 0xe0a4 */
            {8'h00}, /* 0xe0a3 */
            {8'h00}, /* 0xe0a2 */
            {8'h00}, /* 0xe0a1 */
            {8'h00}, /* 0xe0a0 */
            {8'h00}, /* 0xe09f */
            {8'h00}, /* 0xe09e */
            {8'h00}, /* 0xe09d */
            {8'h00}, /* 0xe09c */
            {8'h00}, /* 0xe09b */
            {8'h00}, /* 0xe09a */
            {8'h00}, /* 0xe099 */
            {8'h00}, /* 0xe098 */
            {8'h00}, /* 0xe097 */
            {8'h00}, /* 0xe096 */
            {8'h00}, /* 0xe095 */
            {8'h00}, /* 0xe094 */
            {8'h00}, /* 0xe093 */
            {8'h00}, /* 0xe092 */
            {8'h00}, /* 0xe091 */
            {8'h00}, /* 0xe090 */
            {8'h00}, /* 0xe08f */
            {8'h00}, /* 0xe08e */
            {8'h00}, /* 0xe08d */
            {8'h00}, /* 0xe08c */
            {8'h00}, /* 0xe08b */
            {8'h00}, /* 0xe08a */
            {8'h00}, /* 0xe089 */
            {8'h00}, /* 0xe088 */
            {8'h00}, /* 0xe087 */
            {8'h00}, /* 0xe086 */
            {8'h00}, /* 0xe085 */
            {8'h00}, /* 0xe084 */
            {8'h00}, /* 0xe083 */
            {8'h00}, /* 0xe082 */
            {8'h00}, /* 0xe081 */
            {8'h00}, /* 0xe080 */
            {8'h00}, /* 0xe07f */
            {8'h00}, /* 0xe07e */
            {8'h00}, /* 0xe07d */
            {8'h00}, /* 0xe07c */
            {8'h00}, /* 0xe07b */
            {8'h00}, /* 0xe07a */
            {8'h00}, /* 0xe079 */
            {8'h00}, /* 0xe078 */
            {8'h00}, /* 0xe077 */
            {8'h00}, /* 0xe076 */
            {8'h00}, /* 0xe075 */
            {8'h00}, /* 0xe074 */
            {8'h00}, /* 0xe073 */
            {8'h00}, /* 0xe072 */
            {8'h00}, /* 0xe071 */
            {8'h00}, /* 0xe070 */
            {8'h00}, /* 0xe06f */
            {8'h00}, /* 0xe06e */
            {8'h00}, /* 0xe06d */
            {8'h00}, /* 0xe06c */
            {8'h00}, /* 0xe06b */
            {8'h00}, /* 0xe06a */
            {8'h00}, /* 0xe069 */
            {8'h00}, /* 0xe068 */
            {8'h00}, /* 0xe067 */
            {8'h00}, /* 0xe066 */
            {8'h00}, /* 0xe065 */
            {8'h00}, /* 0xe064 */
            {8'h00}, /* 0xe063 */
            {8'h00}, /* 0xe062 */
            {8'h00}, /* 0xe061 */
            {8'h00}, /* 0xe060 */
            {8'h00}, /* 0xe05f */
            {8'h00}, /* 0xe05e */
            {8'h00}, /* 0xe05d */
            {8'h00}, /* 0xe05c */
            {8'h00}, /* 0xe05b */
            {8'h00}, /* 0xe05a */
            {8'h00}, /* 0xe059 */
            {8'h00}, /* 0xe058 */
            {8'h00}, /* 0xe057 */
            {8'h00}, /* 0xe056 */
            {8'h00}, /* 0xe055 */
            {8'h00}, /* 0xe054 */
            {8'h00}, /* 0xe053 */
            {8'h00}, /* 0xe052 */
            {8'h00}, /* 0xe051 */
            {8'h00}, /* 0xe050 */
            {8'h00}, /* 0xe04f */
            {8'h00}, /* 0xe04e */
            {8'h00}, /* 0xe04d */
            {8'h00}, /* 0xe04c */
            {8'h00}, /* 0xe04b */
            {8'h00}, /* 0xe04a */
            {8'h00}, /* 0xe049 */
            {8'h00}, /* 0xe048 */
            {8'h00}, /* 0xe047 */
            {8'h00}, /* 0xe046 */
            {8'h00}, /* 0xe045 */
            {8'h00}, /* 0xe044 */
            {8'h00}, /* 0xe043 */
            {8'h00}, /* 0xe042 */
            {8'h00}, /* 0xe041 */
            {8'h00}, /* 0xe040 */
            {8'h00}, /* 0xe03f */
            {8'h00}, /* 0xe03e */
            {8'h00}, /* 0xe03d */
            {8'h00}, /* 0xe03c */
            {8'h00}, /* 0xe03b */
            {8'h00}, /* 0xe03a */
            {8'h00}, /* 0xe039 */
            {8'h00}, /* 0xe038 */
            {8'h00}, /* 0xe037 */
            {8'h00}, /* 0xe036 */
            {8'h00}, /* 0xe035 */
            {8'h00}, /* 0xe034 */
            {8'h00}, /* 0xe033 */
            {8'h00}, /* 0xe032 */
            {8'h00}, /* 0xe031 */
            {8'h00}, /* 0xe030 */
            {8'h00}, /* 0xe02f */
            {8'h00}, /* 0xe02e */
            {8'h00}, /* 0xe02d */
            {8'h00}, /* 0xe02c */
            {8'h00}, /* 0xe02b */
            {8'h00}, /* 0xe02a */
            {8'h00}, /* 0xe029 */
            {8'h00}, /* 0xe028 */
            {8'h00}, /* 0xe027 */
            {8'h00}, /* 0xe026 */
            {8'h00}, /* 0xe025 */
            {8'h00}, /* 0xe024 */
            {8'h00}, /* 0xe023 */
            {8'h00}, /* 0xe022 */
            {8'h00}, /* 0xe021 */
            {8'h00}, /* 0xe020 */
            {8'h00}, /* 0xe01f */
            {8'h00}, /* 0xe01e */
            {8'h00}, /* 0xe01d */
            {8'h00}, /* 0xe01c */
            {8'h00}, /* 0xe01b */
            {8'h00}, /* 0xe01a */
            {8'h00}, /* 0xe019 */
            {8'h00}, /* 0xe018 */
            {8'h00}, /* 0xe017 */
            {8'h00}, /* 0xe016 */
            {8'h00}, /* 0xe015 */
            {8'h00}, /* 0xe014 */
            {8'h00}, /* 0xe013 */
            {8'h00}, /* 0xe012 */
            {8'h00}, /* 0xe011 */
            {8'h00}, /* 0xe010 */
            {8'h00}, /* 0xe00f */
            {8'h00}, /* 0xe00e */
            {8'h00}, /* 0xe00d */
            {8'h00}, /* 0xe00c */
            {8'h00}, /* 0xe00b */
            {8'h00}, /* 0xe00a */
            {8'h00}, /* 0xe009 */
            {8'h00}, /* 0xe008 */
            {8'h00}, /* 0xe007 */
            {8'h00}, /* 0xe006 */
            {8'h00}, /* 0xe005 */
            {8'h00}, /* 0xe004 */
            {8'h00}, /* 0xe003 */
            {8'h00}, /* 0xe002 */
            {8'h00}, /* 0xe001 */
            {8'h00}, /* 0xe000 */
            {8'h00}, /* 0xdfff */
            {8'h00}, /* 0xdffe */
            {8'h00}, /* 0xdffd */
            {8'h00}, /* 0xdffc */
            {8'h00}, /* 0xdffb */
            {8'h00}, /* 0xdffa */
            {8'h00}, /* 0xdff9 */
            {8'h00}, /* 0xdff8 */
            {8'h00}, /* 0xdff7 */
            {8'h00}, /* 0xdff6 */
            {8'h00}, /* 0xdff5 */
            {8'h00}, /* 0xdff4 */
            {8'h00}, /* 0xdff3 */
            {8'h00}, /* 0xdff2 */
            {8'h00}, /* 0xdff1 */
            {8'h00}, /* 0xdff0 */
            {8'h00}, /* 0xdfef */
            {8'h00}, /* 0xdfee */
            {8'h00}, /* 0xdfed */
            {8'h00}, /* 0xdfec */
            {8'h00}, /* 0xdfeb */
            {8'h00}, /* 0xdfea */
            {8'h00}, /* 0xdfe9 */
            {8'h00}, /* 0xdfe8 */
            {8'h00}, /* 0xdfe7 */
            {8'h00}, /* 0xdfe6 */
            {8'h00}, /* 0xdfe5 */
            {8'h00}, /* 0xdfe4 */
            {8'h00}, /* 0xdfe3 */
            {8'h00}, /* 0xdfe2 */
            {8'h00}, /* 0xdfe1 */
            {8'h00}, /* 0xdfe0 */
            {8'h00}, /* 0xdfdf */
            {8'h00}, /* 0xdfde */
            {8'h00}, /* 0xdfdd */
            {8'h00}, /* 0xdfdc */
            {8'h00}, /* 0xdfdb */
            {8'h00}, /* 0xdfda */
            {8'h00}, /* 0xdfd9 */
            {8'h00}, /* 0xdfd8 */
            {8'h00}, /* 0xdfd7 */
            {8'h00}, /* 0xdfd6 */
            {8'h00}, /* 0xdfd5 */
            {8'h00}, /* 0xdfd4 */
            {8'h00}, /* 0xdfd3 */
            {8'h00}, /* 0xdfd2 */
            {8'h00}, /* 0xdfd1 */
            {8'h00}, /* 0xdfd0 */
            {8'h00}, /* 0xdfcf */
            {8'h00}, /* 0xdfce */
            {8'h00}, /* 0xdfcd */
            {8'h00}, /* 0xdfcc */
            {8'h00}, /* 0xdfcb */
            {8'h00}, /* 0xdfca */
            {8'h00}, /* 0xdfc9 */
            {8'h00}, /* 0xdfc8 */
            {8'h00}, /* 0xdfc7 */
            {8'h00}, /* 0xdfc6 */
            {8'h00}, /* 0xdfc5 */
            {8'h00}, /* 0xdfc4 */
            {8'h00}, /* 0xdfc3 */
            {8'h00}, /* 0xdfc2 */
            {8'h00}, /* 0xdfc1 */
            {8'h00}, /* 0xdfc0 */
            {8'h00}, /* 0xdfbf */
            {8'h00}, /* 0xdfbe */
            {8'h00}, /* 0xdfbd */
            {8'h00}, /* 0xdfbc */
            {8'h00}, /* 0xdfbb */
            {8'h00}, /* 0xdfba */
            {8'h00}, /* 0xdfb9 */
            {8'h00}, /* 0xdfb8 */
            {8'h00}, /* 0xdfb7 */
            {8'h00}, /* 0xdfb6 */
            {8'h00}, /* 0xdfb5 */
            {8'h00}, /* 0xdfb4 */
            {8'h00}, /* 0xdfb3 */
            {8'h00}, /* 0xdfb2 */
            {8'h00}, /* 0xdfb1 */
            {8'h00}, /* 0xdfb0 */
            {8'h00}, /* 0xdfaf */
            {8'h00}, /* 0xdfae */
            {8'h00}, /* 0xdfad */
            {8'h00}, /* 0xdfac */
            {8'h00}, /* 0xdfab */
            {8'h00}, /* 0xdfaa */
            {8'h00}, /* 0xdfa9 */
            {8'h00}, /* 0xdfa8 */
            {8'h00}, /* 0xdfa7 */
            {8'h00}, /* 0xdfa6 */
            {8'h00}, /* 0xdfa5 */
            {8'h00}, /* 0xdfa4 */
            {8'h00}, /* 0xdfa3 */
            {8'h00}, /* 0xdfa2 */
            {8'h00}, /* 0xdfa1 */
            {8'h00}, /* 0xdfa0 */
            {8'h00}, /* 0xdf9f */
            {8'h00}, /* 0xdf9e */
            {8'h00}, /* 0xdf9d */
            {8'h00}, /* 0xdf9c */
            {8'h00}, /* 0xdf9b */
            {8'h00}, /* 0xdf9a */
            {8'h00}, /* 0xdf99 */
            {8'h00}, /* 0xdf98 */
            {8'h00}, /* 0xdf97 */
            {8'h00}, /* 0xdf96 */
            {8'h00}, /* 0xdf95 */
            {8'h00}, /* 0xdf94 */
            {8'h00}, /* 0xdf93 */
            {8'h00}, /* 0xdf92 */
            {8'h00}, /* 0xdf91 */
            {8'h00}, /* 0xdf90 */
            {8'h00}, /* 0xdf8f */
            {8'h00}, /* 0xdf8e */
            {8'h00}, /* 0xdf8d */
            {8'h00}, /* 0xdf8c */
            {8'h00}, /* 0xdf8b */
            {8'h00}, /* 0xdf8a */
            {8'h00}, /* 0xdf89 */
            {8'h00}, /* 0xdf88 */
            {8'h00}, /* 0xdf87 */
            {8'h00}, /* 0xdf86 */
            {8'h00}, /* 0xdf85 */
            {8'h00}, /* 0xdf84 */
            {8'h00}, /* 0xdf83 */
            {8'h00}, /* 0xdf82 */
            {8'h00}, /* 0xdf81 */
            {8'h00}, /* 0xdf80 */
            {8'h00}, /* 0xdf7f */
            {8'h00}, /* 0xdf7e */
            {8'h00}, /* 0xdf7d */
            {8'h00}, /* 0xdf7c */
            {8'h00}, /* 0xdf7b */
            {8'h00}, /* 0xdf7a */
            {8'h00}, /* 0xdf79 */
            {8'h00}, /* 0xdf78 */
            {8'h00}, /* 0xdf77 */
            {8'h00}, /* 0xdf76 */
            {8'h00}, /* 0xdf75 */
            {8'h00}, /* 0xdf74 */
            {8'h00}, /* 0xdf73 */
            {8'h00}, /* 0xdf72 */
            {8'h00}, /* 0xdf71 */
            {8'h00}, /* 0xdf70 */
            {8'h00}, /* 0xdf6f */
            {8'h00}, /* 0xdf6e */
            {8'h00}, /* 0xdf6d */
            {8'h00}, /* 0xdf6c */
            {8'h00}, /* 0xdf6b */
            {8'h00}, /* 0xdf6a */
            {8'h00}, /* 0xdf69 */
            {8'h00}, /* 0xdf68 */
            {8'h00}, /* 0xdf67 */
            {8'h00}, /* 0xdf66 */
            {8'h00}, /* 0xdf65 */
            {8'h00}, /* 0xdf64 */
            {8'h00}, /* 0xdf63 */
            {8'h00}, /* 0xdf62 */
            {8'h00}, /* 0xdf61 */
            {8'h00}, /* 0xdf60 */
            {8'h00}, /* 0xdf5f */
            {8'h00}, /* 0xdf5e */
            {8'h00}, /* 0xdf5d */
            {8'h00}, /* 0xdf5c */
            {8'h00}, /* 0xdf5b */
            {8'h00}, /* 0xdf5a */
            {8'h00}, /* 0xdf59 */
            {8'h00}, /* 0xdf58 */
            {8'h00}, /* 0xdf57 */
            {8'h00}, /* 0xdf56 */
            {8'h00}, /* 0xdf55 */
            {8'h00}, /* 0xdf54 */
            {8'h00}, /* 0xdf53 */
            {8'h00}, /* 0xdf52 */
            {8'h00}, /* 0xdf51 */
            {8'h00}, /* 0xdf50 */
            {8'h00}, /* 0xdf4f */
            {8'h00}, /* 0xdf4e */
            {8'h00}, /* 0xdf4d */
            {8'h00}, /* 0xdf4c */
            {8'h00}, /* 0xdf4b */
            {8'h00}, /* 0xdf4a */
            {8'h00}, /* 0xdf49 */
            {8'h00}, /* 0xdf48 */
            {8'h00}, /* 0xdf47 */
            {8'h00}, /* 0xdf46 */
            {8'h00}, /* 0xdf45 */
            {8'h00}, /* 0xdf44 */
            {8'h00}, /* 0xdf43 */
            {8'h00}, /* 0xdf42 */
            {8'h00}, /* 0xdf41 */
            {8'h00}, /* 0xdf40 */
            {8'h00}, /* 0xdf3f */
            {8'h00}, /* 0xdf3e */
            {8'h00}, /* 0xdf3d */
            {8'h00}, /* 0xdf3c */
            {8'h00}, /* 0xdf3b */
            {8'h00}, /* 0xdf3a */
            {8'h00}, /* 0xdf39 */
            {8'h00}, /* 0xdf38 */
            {8'h00}, /* 0xdf37 */
            {8'h00}, /* 0xdf36 */
            {8'h00}, /* 0xdf35 */
            {8'h00}, /* 0xdf34 */
            {8'h00}, /* 0xdf33 */
            {8'h00}, /* 0xdf32 */
            {8'h00}, /* 0xdf31 */
            {8'h00}, /* 0xdf30 */
            {8'h00}, /* 0xdf2f */
            {8'h00}, /* 0xdf2e */
            {8'h00}, /* 0xdf2d */
            {8'h00}, /* 0xdf2c */
            {8'h00}, /* 0xdf2b */
            {8'h00}, /* 0xdf2a */
            {8'h00}, /* 0xdf29 */
            {8'h00}, /* 0xdf28 */
            {8'h00}, /* 0xdf27 */
            {8'h00}, /* 0xdf26 */
            {8'h00}, /* 0xdf25 */
            {8'h00}, /* 0xdf24 */
            {8'h00}, /* 0xdf23 */
            {8'h00}, /* 0xdf22 */
            {8'h00}, /* 0xdf21 */
            {8'h00}, /* 0xdf20 */
            {8'h00}, /* 0xdf1f */
            {8'h00}, /* 0xdf1e */
            {8'h00}, /* 0xdf1d */
            {8'h00}, /* 0xdf1c */
            {8'h00}, /* 0xdf1b */
            {8'h00}, /* 0xdf1a */
            {8'h00}, /* 0xdf19 */
            {8'h00}, /* 0xdf18 */
            {8'h00}, /* 0xdf17 */
            {8'h00}, /* 0xdf16 */
            {8'h00}, /* 0xdf15 */
            {8'h00}, /* 0xdf14 */
            {8'h00}, /* 0xdf13 */
            {8'h00}, /* 0xdf12 */
            {8'h00}, /* 0xdf11 */
            {8'h00}, /* 0xdf10 */
            {8'h00}, /* 0xdf0f */
            {8'h00}, /* 0xdf0e */
            {8'h00}, /* 0xdf0d */
            {8'h00}, /* 0xdf0c */
            {8'h00}, /* 0xdf0b */
            {8'h00}, /* 0xdf0a */
            {8'h00}, /* 0xdf09 */
            {8'h00}, /* 0xdf08 */
            {8'h00}, /* 0xdf07 */
            {8'h00}, /* 0xdf06 */
            {8'h00}, /* 0xdf05 */
            {8'h00}, /* 0xdf04 */
            {8'h00}, /* 0xdf03 */
            {8'h00}, /* 0xdf02 */
            {8'h00}, /* 0xdf01 */
            {8'h00}, /* 0xdf00 */
            {8'h00}, /* 0xdeff */
            {8'h00}, /* 0xdefe */
            {8'h00}, /* 0xdefd */
            {8'h00}, /* 0xdefc */
            {8'h00}, /* 0xdefb */
            {8'h00}, /* 0xdefa */
            {8'h00}, /* 0xdef9 */
            {8'h00}, /* 0xdef8 */
            {8'h00}, /* 0xdef7 */
            {8'h00}, /* 0xdef6 */
            {8'h00}, /* 0xdef5 */
            {8'h00}, /* 0xdef4 */
            {8'h00}, /* 0xdef3 */
            {8'h00}, /* 0xdef2 */
            {8'h00}, /* 0xdef1 */
            {8'h00}, /* 0xdef0 */
            {8'h00}, /* 0xdeef */
            {8'h00}, /* 0xdeee */
            {8'h00}, /* 0xdeed */
            {8'h00}, /* 0xdeec */
            {8'h00}, /* 0xdeeb */
            {8'h00}, /* 0xdeea */
            {8'h00}, /* 0xdee9 */
            {8'h00}, /* 0xdee8 */
            {8'h00}, /* 0xdee7 */
            {8'h00}, /* 0xdee6 */
            {8'h00}, /* 0xdee5 */
            {8'h00}, /* 0xdee4 */
            {8'h00}, /* 0xdee3 */
            {8'h00}, /* 0xdee2 */
            {8'h00}, /* 0xdee1 */
            {8'h00}, /* 0xdee0 */
            {8'h00}, /* 0xdedf */
            {8'h00}, /* 0xdede */
            {8'h00}, /* 0xdedd */
            {8'h00}, /* 0xdedc */
            {8'h00}, /* 0xdedb */
            {8'h00}, /* 0xdeda */
            {8'h00}, /* 0xded9 */
            {8'h00}, /* 0xded8 */
            {8'h00}, /* 0xded7 */
            {8'h00}, /* 0xded6 */
            {8'h00}, /* 0xded5 */
            {8'h00}, /* 0xded4 */
            {8'h00}, /* 0xded3 */
            {8'h00}, /* 0xded2 */
            {8'h00}, /* 0xded1 */
            {8'h00}, /* 0xded0 */
            {8'h00}, /* 0xdecf */
            {8'h00}, /* 0xdece */
            {8'h00}, /* 0xdecd */
            {8'h00}, /* 0xdecc */
            {8'h00}, /* 0xdecb */
            {8'h00}, /* 0xdeca */
            {8'h00}, /* 0xdec9 */
            {8'h00}, /* 0xdec8 */
            {8'h00}, /* 0xdec7 */
            {8'h00}, /* 0xdec6 */
            {8'h00}, /* 0xdec5 */
            {8'h00}, /* 0xdec4 */
            {8'h00}, /* 0xdec3 */
            {8'h00}, /* 0xdec2 */
            {8'h00}, /* 0xdec1 */
            {8'h00}, /* 0xdec0 */
            {8'h00}, /* 0xdebf */
            {8'h00}, /* 0xdebe */
            {8'h00}, /* 0xdebd */
            {8'h00}, /* 0xdebc */
            {8'h00}, /* 0xdebb */
            {8'h00}, /* 0xdeba */
            {8'h00}, /* 0xdeb9 */
            {8'h00}, /* 0xdeb8 */
            {8'h00}, /* 0xdeb7 */
            {8'h00}, /* 0xdeb6 */
            {8'h00}, /* 0xdeb5 */
            {8'h00}, /* 0xdeb4 */
            {8'h00}, /* 0xdeb3 */
            {8'h00}, /* 0xdeb2 */
            {8'h00}, /* 0xdeb1 */
            {8'h00}, /* 0xdeb0 */
            {8'h00}, /* 0xdeaf */
            {8'h00}, /* 0xdeae */
            {8'h00}, /* 0xdead */
            {8'h00}, /* 0xdeac */
            {8'h00}, /* 0xdeab */
            {8'h00}, /* 0xdeaa */
            {8'h00}, /* 0xdea9 */
            {8'h00}, /* 0xdea8 */
            {8'h00}, /* 0xdea7 */
            {8'h00}, /* 0xdea6 */
            {8'h00}, /* 0xdea5 */
            {8'h00}, /* 0xdea4 */
            {8'h00}, /* 0xdea3 */
            {8'h00}, /* 0xdea2 */
            {8'h00}, /* 0xdea1 */
            {8'h00}, /* 0xdea0 */
            {8'h00}, /* 0xde9f */
            {8'h00}, /* 0xde9e */
            {8'h00}, /* 0xde9d */
            {8'h00}, /* 0xde9c */
            {8'h00}, /* 0xde9b */
            {8'h00}, /* 0xde9a */
            {8'h00}, /* 0xde99 */
            {8'h00}, /* 0xde98 */
            {8'h00}, /* 0xde97 */
            {8'h00}, /* 0xde96 */
            {8'h00}, /* 0xde95 */
            {8'h00}, /* 0xde94 */
            {8'h00}, /* 0xde93 */
            {8'h00}, /* 0xde92 */
            {8'h00}, /* 0xde91 */
            {8'h00}, /* 0xde90 */
            {8'h00}, /* 0xde8f */
            {8'h00}, /* 0xde8e */
            {8'h00}, /* 0xde8d */
            {8'h00}, /* 0xde8c */
            {8'h00}, /* 0xde8b */
            {8'h00}, /* 0xde8a */
            {8'h00}, /* 0xde89 */
            {8'h00}, /* 0xde88 */
            {8'h00}, /* 0xde87 */
            {8'h00}, /* 0xde86 */
            {8'h00}, /* 0xde85 */
            {8'h00}, /* 0xde84 */
            {8'h00}, /* 0xde83 */
            {8'h00}, /* 0xde82 */
            {8'h00}, /* 0xde81 */
            {8'h00}, /* 0xde80 */
            {8'h00}, /* 0xde7f */
            {8'h00}, /* 0xde7e */
            {8'h00}, /* 0xde7d */
            {8'h00}, /* 0xde7c */
            {8'h00}, /* 0xde7b */
            {8'h00}, /* 0xde7a */
            {8'h00}, /* 0xde79 */
            {8'h00}, /* 0xde78 */
            {8'h00}, /* 0xde77 */
            {8'h00}, /* 0xde76 */
            {8'h00}, /* 0xde75 */
            {8'h00}, /* 0xde74 */
            {8'h00}, /* 0xde73 */
            {8'h00}, /* 0xde72 */
            {8'h00}, /* 0xde71 */
            {8'h00}, /* 0xde70 */
            {8'h00}, /* 0xde6f */
            {8'h00}, /* 0xde6e */
            {8'h00}, /* 0xde6d */
            {8'h00}, /* 0xde6c */
            {8'h00}, /* 0xde6b */
            {8'h00}, /* 0xde6a */
            {8'h00}, /* 0xde69 */
            {8'h00}, /* 0xde68 */
            {8'h00}, /* 0xde67 */
            {8'h00}, /* 0xde66 */
            {8'h00}, /* 0xde65 */
            {8'h00}, /* 0xde64 */
            {8'h00}, /* 0xde63 */
            {8'h00}, /* 0xde62 */
            {8'h00}, /* 0xde61 */
            {8'h00}, /* 0xde60 */
            {8'h00}, /* 0xde5f */
            {8'h00}, /* 0xde5e */
            {8'h00}, /* 0xde5d */
            {8'h00}, /* 0xde5c */
            {8'h00}, /* 0xde5b */
            {8'h00}, /* 0xde5a */
            {8'h00}, /* 0xde59 */
            {8'h00}, /* 0xde58 */
            {8'h00}, /* 0xde57 */
            {8'h00}, /* 0xde56 */
            {8'h00}, /* 0xde55 */
            {8'h00}, /* 0xde54 */
            {8'h00}, /* 0xde53 */
            {8'h00}, /* 0xde52 */
            {8'h00}, /* 0xde51 */
            {8'h00}, /* 0xde50 */
            {8'h00}, /* 0xde4f */
            {8'h00}, /* 0xde4e */
            {8'h00}, /* 0xde4d */
            {8'h00}, /* 0xde4c */
            {8'h00}, /* 0xde4b */
            {8'h00}, /* 0xde4a */
            {8'h00}, /* 0xde49 */
            {8'h00}, /* 0xde48 */
            {8'h00}, /* 0xde47 */
            {8'h00}, /* 0xde46 */
            {8'h00}, /* 0xde45 */
            {8'h00}, /* 0xde44 */
            {8'h00}, /* 0xde43 */
            {8'h00}, /* 0xde42 */
            {8'h00}, /* 0xde41 */
            {8'h00}, /* 0xde40 */
            {8'h00}, /* 0xde3f */
            {8'h00}, /* 0xde3e */
            {8'h00}, /* 0xde3d */
            {8'h00}, /* 0xde3c */
            {8'h00}, /* 0xde3b */
            {8'h00}, /* 0xde3a */
            {8'h00}, /* 0xde39 */
            {8'h00}, /* 0xde38 */
            {8'h00}, /* 0xde37 */
            {8'h00}, /* 0xde36 */
            {8'h00}, /* 0xde35 */
            {8'h00}, /* 0xde34 */
            {8'h00}, /* 0xde33 */
            {8'h00}, /* 0xde32 */
            {8'h00}, /* 0xde31 */
            {8'h00}, /* 0xde30 */
            {8'h00}, /* 0xde2f */
            {8'h00}, /* 0xde2e */
            {8'h00}, /* 0xde2d */
            {8'h00}, /* 0xde2c */
            {8'h00}, /* 0xde2b */
            {8'h00}, /* 0xde2a */
            {8'h00}, /* 0xde29 */
            {8'h00}, /* 0xde28 */
            {8'h00}, /* 0xde27 */
            {8'h00}, /* 0xde26 */
            {8'h00}, /* 0xde25 */
            {8'h00}, /* 0xde24 */
            {8'h00}, /* 0xde23 */
            {8'h00}, /* 0xde22 */
            {8'h00}, /* 0xde21 */
            {8'h00}, /* 0xde20 */
            {8'h00}, /* 0xde1f */
            {8'h00}, /* 0xde1e */
            {8'h00}, /* 0xde1d */
            {8'h00}, /* 0xde1c */
            {8'h00}, /* 0xde1b */
            {8'h00}, /* 0xde1a */
            {8'h00}, /* 0xde19 */
            {8'h00}, /* 0xde18 */
            {8'h00}, /* 0xde17 */
            {8'h00}, /* 0xde16 */
            {8'h00}, /* 0xde15 */
            {8'h00}, /* 0xde14 */
            {8'h00}, /* 0xde13 */
            {8'h00}, /* 0xde12 */
            {8'h00}, /* 0xde11 */
            {8'h00}, /* 0xde10 */
            {8'h00}, /* 0xde0f */
            {8'h00}, /* 0xde0e */
            {8'h00}, /* 0xde0d */
            {8'h00}, /* 0xde0c */
            {8'h00}, /* 0xde0b */
            {8'h00}, /* 0xde0a */
            {8'h00}, /* 0xde09 */
            {8'h00}, /* 0xde08 */
            {8'h00}, /* 0xde07 */
            {8'h00}, /* 0xde06 */
            {8'h00}, /* 0xde05 */
            {8'h00}, /* 0xde04 */
            {8'h00}, /* 0xde03 */
            {8'h00}, /* 0xde02 */
            {8'h00}, /* 0xde01 */
            {8'h00}, /* 0xde00 */
            {8'h00}, /* 0xddff */
            {8'h00}, /* 0xddfe */
            {8'h00}, /* 0xddfd */
            {8'h00}, /* 0xddfc */
            {8'h00}, /* 0xddfb */
            {8'h00}, /* 0xddfa */
            {8'h00}, /* 0xddf9 */
            {8'h00}, /* 0xddf8 */
            {8'h00}, /* 0xddf7 */
            {8'h00}, /* 0xddf6 */
            {8'h00}, /* 0xddf5 */
            {8'h00}, /* 0xddf4 */
            {8'h00}, /* 0xddf3 */
            {8'h00}, /* 0xddf2 */
            {8'h00}, /* 0xddf1 */
            {8'h00}, /* 0xddf0 */
            {8'h00}, /* 0xddef */
            {8'h00}, /* 0xddee */
            {8'h00}, /* 0xdded */
            {8'h00}, /* 0xddec */
            {8'h00}, /* 0xddeb */
            {8'h00}, /* 0xddea */
            {8'h00}, /* 0xdde9 */
            {8'h00}, /* 0xdde8 */
            {8'h00}, /* 0xdde7 */
            {8'h00}, /* 0xdde6 */
            {8'h00}, /* 0xdde5 */
            {8'h00}, /* 0xdde4 */
            {8'h00}, /* 0xdde3 */
            {8'h00}, /* 0xdde2 */
            {8'h00}, /* 0xdde1 */
            {8'h00}, /* 0xdde0 */
            {8'h00}, /* 0xdddf */
            {8'h00}, /* 0xddde */
            {8'h00}, /* 0xdddd */
            {8'h00}, /* 0xdddc */
            {8'h00}, /* 0xdddb */
            {8'h00}, /* 0xddda */
            {8'h00}, /* 0xddd9 */
            {8'h00}, /* 0xddd8 */
            {8'h00}, /* 0xddd7 */
            {8'h00}, /* 0xddd6 */
            {8'h00}, /* 0xddd5 */
            {8'h00}, /* 0xddd4 */
            {8'h00}, /* 0xddd3 */
            {8'h00}, /* 0xddd2 */
            {8'h00}, /* 0xddd1 */
            {8'h00}, /* 0xddd0 */
            {8'h00}, /* 0xddcf */
            {8'h00}, /* 0xddce */
            {8'h00}, /* 0xddcd */
            {8'h00}, /* 0xddcc */
            {8'h00}, /* 0xddcb */
            {8'h00}, /* 0xddca */
            {8'h00}, /* 0xddc9 */
            {8'h00}, /* 0xddc8 */
            {8'h00}, /* 0xddc7 */
            {8'h00}, /* 0xddc6 */
            {8'h00}, /* 0xddc5 */
            {8'h00}, /* 0xddc4 */
            {8'h00}, /* 0xddc3 */
            {8'h00}, /* 0xddc2 */
            {8'h00}, /* 0xddc1 */
            {8'h00}, /* 0xddc0 */
            {8'h00}, /* 0xddbf */
            {8'h00}, /* 0xddbe */
            {8'h00}, /* 0xddbd */
            {8'h00}, /* 0xddbc */
            {8'h00}, /* 0xddbb */
            {8'h00}, /* 0xddba */
            {8'h00}, /* 0xddb9 */
            {8'h00}, /* 0xddb8 */
            {8'h00}, /* 0xddb7 */
            {8'h00}, /* 0xddb6 */
            {8'h00}, /* 0xddb5 */
            {8'h00}, /* 0xddb4 */
            {8'h00}, /* 0xddb3 */
            {8'h00}, /* 0xddb2 */
            {8'h00}, /* 0xddb1 */
            {8'h00}, /* 0xddb0 */
            {8'h00}, /* 0xddaf */
            {8'h00}, /* 0xddae */
            {8'h00}, /* 0xddad */
            {8'h00}, /* 0xddac */
            {8'h00}, /* 0xddab */
            {8'h00}, /* 0xddaa */
            {8'h00}, /* 0xdda9 */
            {8'h00}, /* 0xdda8 */
            {8'h00}, /* 0xdda7 */
            {8'h00}, /* 0xdda6 */
            {8'h00}, /* 0xdda5 */
            {8'h00}, /* 0xdda4 */
            {8'h00}, /* 0xdda3 */
            {8'h00}, /* 0xdda2 */
            {8'h00}, /* 0xdda1 */
            {8'h00}, /* 0xdda0 */
            {8'h00}, /* 0xdd9f */
            {8'h00}, /* 0xdd9e */
            {8'h00}, /* 0xdd9d */
            {8'h00}, /* 0xdd9c */
            {8'h00}, /* 0xdd9b */
            {8'h00}, /* 0xdd9a */
            {8'h00}, /* 0xdd99 */
            {8'h00}, /* 0xdd98 */
            {8'h00}, /* 0xdd97 */
            {8'h00}, /* 0xdd96 */
            {8'h00}, /* 0xdd95 */
            {8'h00}, /* 0xdd94 */
            {8'h00}, /* 0xdd93 */
            {8'h00}, /* 0xdd92 */
            {8'h00}, /* 0xdd91 */
            {8'h00}, /* 0xdd90 */
            {8'h00}, /* 0xdd8f */
            {8'h00}, /* 0xdd8e */
            {8'h00}, /* 0xdd8d */
            {8'h00}, /* 0xdd8c */
            {8'h00}, /* 0xdd8b */
            {8'h00}, /* 0xdd8a */
            {8'h00}, /* 0xdd89 */
            {8'h00}, /* 0xdd88 */
            {8'h00}, /* 0xdd87 */
            {8'h00}, /* 0xdd86 */
            {8'h00}, /* 0xdd85 */
            {8'h00}, /* 0xdd84 */
            {8'h00}, /* 0xdd83 */
            {8'h00}, /* 0xdd82 */
            {8'h00}, /* 0xdd81 */
            {8'h00}, /* 0xdd80 */
            {8'h00}, /* 0xdd7f */
            {8'h00}, /* 0xdd7e */
            {8'h00}, /* 0xdd7d */
            {8'h00}, /* 0xdd7c */
            {8'h00}, /* 0xdd7b */
            {8'h00}, /* 0xdd7a */
            {8'h00}, /* 0xdd79 */
            {8'h00}, /* 0xdd78 */
            {8'h00}, /* 0xdd77 */
            {8'h00}, /* 0xdd76 */
            {8'h00}, /* 0xdd75 */
            {8'h00}, /* 0xdd74 */
            {8'h00}, /* 0xdd73 */
            {8'h00}, /* 0xdd72 */
            {8'h00}, /* 0xdd71 */
            {8'h00}, /* 0xdd70 */
            {8'h00}, /* 0xdd6f */
            {8'h00}, /* 0xdd6e */
            {8'h00}, /* 0xdd6d */
            {8'h00}, /* 0xdd6c */
            {8'h00}, /* 0xdd6b */
            {8'h00}, /* 0xdd6a */
            {8'h00}, /* 0xdd69 */
            {8'h00}, /* 0xdd68 */
            {8'h00}, /* 0xdd67 */
            {8'h00}, /* 0xdd66 */
            {8'h00}, /* 0xdd65 */
            {8'h00}, /* 0xdd64 */
            {8'h00}, /* 0xdd63 */
            {8'h00}, /* 0xdd62 */
            {8'h00}, /* 0xdd61 */
            {8'h00}, /* 0xdd60 */
            {8'h00}, /* 0xdd5f */
            {8'h00}, /* 0xdd5e */
            {8'h00}, /* 0xdd5d */
            {8'h00}, /* 0xdd5c */
            {8'h00}, /* 0xdd5b */
            {8'h00}, /* 0xdd5a */
            {8'h00}, /* 0xdd59 */
            {8'h00}, /* 0xdd58 */
            {8'h00}, /* 0xdd57 */
            {8'h00}, /* 0xdd56 */
            {8'h00}, /* 0xdd55 */
            {8'h00}, /* 0xdd54 */
            {8'h00}, /* 0xdd53 */
            {8'h00}, /* 0xdd52 */
            {8'h00}, /* 0xdd51 */
            {8'h00}, /* 0xdd50 */
            {8'h00}, /* 0xdd4f */
            {8'h00}, /* 0xdd4e */
            {8'h00}, /* 0xdd4d */
            {8'h00}, /* 0xdd4c */
            {8'h00}, /* 0xdd4b */
            {8'h00}, /* 0xdd4a */
            {8'h00}, /* 0xdd49 */
            {8'h00}, /* 0xdd48 */
            {8'h00}, /* 0xdd47 */
            {8'h00}, /* 0xdd46 */
            {8'h00}, /* 0xdd45 */
            {8'h00}, /* 0xdd44 */
            {8'h00}, /* 0xdd43 */
            {8'h00}, /* 0xdd42 */
            {8'h00}, /* 0xdd41 */
            {8'h00}, /* 0xdd40 */
            {8'h00}, /* 0xdd3f */
            {8'h00}, /* 0xdd3e */
            {8'h00}, /* 0xdd3d */
            {8'h00}, /* 0xdd3c */
            {8'h00}, /* 0xdd3b */
            {8'h00}, /* 0xdd3a */
            {8'h00}, /* 0xdd39 */
            {8'h00}, /* 0xdd38 */
            {8'h00}, /* 0xdd37 */
            {8'h00}, /* 0xdd36 */
            {8'h00}, /* 0xdd35 */
            {8'h00}, /* 0xdd34 */
            {8'h00}, /* 0xdd33 */
            {8'h00}, /* 0xdd32 */
            {8'h00}, /* 0xdd31 */
            {8'h00}, /* 0xdd30 */
            {8'h00}, /* 0xdd2f */
            {8'h00}, /* 0xdd2e */
            {8'h00}, /* 0xdd2d */
            {8'h00}, /* 0xdd2c */
            {8'h00}, /* 0xdd2b */
            {8'h00}, /* 0xdd2a */
            {8'h00}, /* 0xdd29 */
            {8'h00}, /* 0xdd28 */
            {8'h00}, /* 0xdd27 */
            {8'h00}, /* 0xdd26 */
            {8'h00}, /* 0xdd25 */
            {8'h00}, /* 0xdd24 */
            {8'h00}, /* 0xdd23 */
            {8'h00}, /* 0xdd22 */
            {8'h00}, /* 0xdd21 */
            {8'h00}, /* 0xdd20 */
            {8'h00}, /* 0xdd1f */
            {8'h00}, /* 0xdd1e */
            {8'h00}, /* 0xdd1d */
            {8'h00}, /* 0xdd1c */
            {8'h00}, /* 0xdd1b */
            {8'h00}, /* 0xdd1a */
            {8'h00}, /* 0xdd19 */
            {8'h00}, /* 0xdd18 */
            {8'h00}, /* 0xdd17 */
            {8'h00}, /* 0xdd16 */
            {8'h00}, /* 0xdd15 */
            {8'h00}, /* 0xdd14 */
            {8'h00}, /* 0xdd13 */
            {8'h00}, /* 0xdd12 */
            {8'h00}, /* 0xdd11 */
            {8'h00}, /* 0xdd10 */
            {8'h00}, /* 0xdd0f */
            {8'h00}, /* 0xdd0e */
            {8'h00}, /* 0xdd0d */
            {8'h00}, /* 0xdd0c */
            {8'h00}, /* 0xdd0b */
            {8'h00}, /* 0xdd0a */
            {8'h00}, /* 0xdd09 */
            {8'h00}, /* 0xdd08 */
            {8'h00}, /* 0xdd07 */
            {8'h00}, /* 0xdd06 */
            {8'h00}, /* 0xdd05 */
            {8'h00}, /* 0xdd04 */
            {8'h00}, /* 0xdd03 */
            {8'h00}, /* 0xdd02 */
            {8'h00}, /* 0xdd01 */
            {8'h00}, /* 0xdd00 */
            {8'h00}, /* 0xdcff */
            {8'h00}, /* 0xdcfe */
            {8'h00}, /* 0xdcfd */
            {8'h00}, /* 0xdcfc */
            {8'h00}, /* 0xdcfb */
            {8'h00}, /* 0xdcfa */
            {8'h00}, /* 0xdcf9 */
            {8'h00}, /* 0xdcf8 */
            {8'h00}, /* 0xdcf7 */
            {8'h00}, /* 0xdcf6 */
            {8'h00}, /* 0xdcf5 */
            {8'h00}, /* 0xdcf4 */
            {8'h00}, /* 0xdcf3 */
            {8'h00}, /* 0xdcf2 */
            {8'h00}, /* 0xdcf1 */
            {8'h00}, /* 0xdcf0 */
            {8'h00}, /* 0xdcef */
            {8'h00}, /* 0xdcee */
            {8'h00}, /* 0xdced */
            {8'h00}, /* 0xdcec */
            {8'h00}, /* 0xdceb */
            {8'h00}, /* 0xdcea */
            {8'h00}, /* 0xdce9 */
            {8'h00}, /* 0xdce8 */
            {8'h00}, /* 0xdce7 */
            {8'h00}, /* 0xdce6 */
            {8'h00}, /* 0xdce5 */
            {8'h00}, /* 0xdce4 */
            {8'h00}, /* 0xdce3 */
            {8'h00}, /* 0xdce2 */
            {8'h00}, /* 0xdce1 */
            {8'h00}, /* 0xdce0 */
            {8'h00}, /* 0xdcdf */
            {8'h00}, /* 0xdcde */
            {8'h00}, /* 0xdcdd */
            {8'h00}, /* 0xdcdc */
            {8'h00}, /* 0xdcdb */
            {8'h00}, /* 0xdcda */
            {8'h00}, /* 0xdcd9 */
            {8'h00}, /* 0xdcd8 */
            {8'h00}, /* 0xdcd7 */
            {8'h00}, /* 0xdcd6 */
            {8'h00}, /* 0xdcd5 */
            {8'h00}, /* 0xdcd4 */
            {8'h00}, /* 0xdcd3 */
            {8'h00}, /* 0xdcd2 */
            {8'h00}, /* 0xdcd1 */
            {8'h00}, /* 0xdcd0 */
            {8'h00}, /* 0xdccf */
            {8'h00}, /* 0xdcce */
            {8'h00}, /* 0xdccd */
            {8'h00}, /* 0xdccc */
            {8'h00}, /* 0xdccb */
            {8'h00}, /* 0xdcca */
            {8'h00}, /* 0xdcc9 */
            {8'h00}, /* 0xdcc8 */
            {8'h00}, /* 0xdcc7 */
            {8'h00}, /* 0xdcc6 */
            {8'h00}, /* 0xdcc5 */
            {8'h00}, /* 0xdcc4 */
            {8'h00}, /* 0xdcc3 */
            {8'h00}, /* 0xdcc2 */
            {8'h00}, /* 0xdcc1 */
            {8'h00}, /* 0xdcc0 */
            {8'h00}, /* 0xdcbf */
            {8'h00}, /* 0xdcbe */
            {8'h00}, /* 0xdcbd */
            {8'h00}, /* 0xdcbc */
            {8'h00}, /* 0xdcbb */
            {8'h00}, /* 0xdcba */
            {8'h00}, /* 0xdcb9 */
            {8'h00}, /* 0xdcb8 */
            {8'h00}, /* 0xdcb7 */
            {8'h00}, /* 0xdcb6 */
            {8'h00}, /* 0xdcb5 */
            {8'h00}, /* 0xdcb4 */
            {8'h00}, /* 0xdcb3 */
            {8'h00}, /* 0xdcb2 */
            {8'h00}, /* 0xdcb1 */
            {8'h00}, /* 0xdcb0 */
            {8'h00}, /* 0xdcaf */
            {8'h00}, /* 0xdcae */
            {8'h00}, /* 0xdcad */
            {8'h00}, /* 0xdcac */
            {8'h00}, /* 0xdcab */
            {8'h00}, /* 0xdcaa */
            {8'h00}, /* 0xdca9 */
            {8'h00}, /* 0xdca8 */
            {8'h00}, /* 0xdca7 */
            {8'h00}, /* 0xdca6 */
            {8'h00}, /* 0xdca5 */
            {8'h00}, /* 0xdca4 */
            {8'h00}, /* 0xdca3 */
            {8'h00}, /* 0xdca2 */
            {8'h00}, /* 0xdca1 */
            {8'h00}, /* 0xdca0 */
            {8'h00}, /* 0xdc9f */
            {8'h00}, /* 0xdc9e */
            {8'h00}, /* 0xdc9d */
            {8'h00}, /* 0xdc9c */
            {8'h00}, /* 0xdc9b */
            {8'h00}, /* 0xdc9a */
            {8'h00}, /* 0xdc99 */
            {8'h00}, /* 0xdc98 */
            {8'h00}, /* 0xdc97 */
            {8'h00}, /* 0xdc96 */
            {8'h00}, /* 0xdc95 */
            {8'h00}, /* 0xdc94 */
            {8'h00}, /* 0xdc93 */
            {8'h00}, /* 0xdc92 */
            {8'h00}, /* 0xdc91 */
            {8'h00}, /* 0xdc90 */
            {8'h00}, /* 0xdc8f */
            {8'h00}, /* 0xdc8e */
            {8'h00}, /* 0xdc8d */
            {8'h00}, /* 0xdc8c */
            {8'h00}, /* 0xdc8b */
            {8'h00}, /* 0xdc8a */
            {8'h00}, /* 0xdc89 */
            {8'h00}, /* 0xdc88 */
            {8'h00}, /* 0xdc87 */
            {8'h00}, /* 0xdc86 */
            {8'h00}, /* 0xdc85 */
            {8'h00}, /* 0xdc84 */
            {8'h00}, /* 0xdc83 */
            {8'h00}, /* 0xdc82 */
            {8'h00}, /* 0xdc81 */
            {8'h00}, /* 0xdc80 */
            {8'h00}, /* 0xdc7f */
            {8'h00}, /* 0xdc7e */
            {8'h00}, /* 0xdc7d */
            {8'h00}, /* 0xdc7c */
            {8'h00}, /* 0xdc7b */
            {8'h00}, /* 0xdc7a */
            {8'h00}, /* 0xdc79 */
            {8'h00}, /* 0xdc78 */
            {8'h00}, /* 0xdc77 */
            {8'h00}, /* 0xdc76 */
            {8'h00}, /* 0xdc75 */
            {8'h00}, /* 0xdc74 */
            {8'h00}, /* 0xdc73 */
            {8'h00}, /* 0xdc72 */
            {8'h00}, /* 0xdc71 */
            {8'h00}, /* 0xdc70 */
            {8'h00}, /* 0xdc6f */
            {8'h00}, /* 0xdc6e */
            {8'h00}, /* 0xdc6d */
            {8'h00}, /* 0xdc6c */
            {8'h00}, /* 0xdc6b */
            {8'h00}, /* 0xdc6a */
            {8'h00}, /* 0xdc69 */
            {8'h00}, /* 0xdc68 */
            {8'h00}, /* 0xdc67 */
            {8'h00}, /* 0xdc66 */
            {8'h00}, /* 0xdc65 */
            {8'h00}, /* 0xdc64 */
            {8'h00}, /* 0xdc63 */
            {8'h00}, /* 0xdc62 */
            {8'h00}, /* 0xdc61 */
            {8'h00}, /* 0xdc60 */
            {8'h00}, /* 0xdc5f */
            {8'h00}, /* 0xdc5e */
            {8'h00}, /* 0xdc5d */
            {8'h00}, /* 0xdc5c */
            {8'h00}, /* 0xdc5b */
            {8'h00}, /* 0xdc5a */
            {8'h00}, /* 0xdc59 */
            {8'h00}, /* 0xdc58 */
            {8'h00}, /* 0xdc57 */
            {8'h00}, /* 0xdc56 */
            {8'h00}, /* 0xdc55 */
            {8'h00}, /* 0xdc54 */
            {8'h00}, /* 0xdc53 */
            {8'h00}, /* 0xdc52 */
            {8'h00}, /* 0xdc51 */
            {8'h00}, /* 0xdc50 */
            {8'h00}, /* 0xdc4f */
            {8'h00}, /* 0xdc4e */
            {8'h00}, /* 0xdc4d */
            {8'h00}, /* 0xdc4c */
            {8'h00}, /* 0xdc4b */
            {8'h00}, /* 0xdc4a */
            {8'h00}, /* 0xdc49 */
            {8'h00}, /* 0xdc48 */
            {8'h00}, /* 0xdc47 */
            {8'h00}, /* 0xdc46 */
            {8'h00}, /* 0xdc45 */
            {8'h00}, /* 0xdc44 */
            {8'h00}, /* 0xdc43 */
            {8'h00}, /* 0xdc42 */
            {8'h00}, /* 0xdc41 */
            {8'h00}, /* 0xdc40 */
            {8'h00}, /* 0xdc3f */
            {8'h00}, /* 0xdc3e */
            {8'h00}, /* 0xdc3d */
            {8'h00}, /* 0xdc3c */
            {8'h00}, /* 0xdc3b */
            {8'h00}, /* 0xdc3a */
            {8'h00}, /* 0xdc39 */
            {8'h00}, /* 0xdc38 */
            {8'h00}, /* 0xdc37 */
            {8'h00}, /* 0xdc36 */
            {8'h00}, /* 0xdc35 */
            {8'h00}, /* 0xdc34 */
            {8'h00}, /* 0xdc33 */
            {8'h00}, /* 0xdc32 */
            {8'h00}, /* 0xdc31 */
            {8'h00}, /* 0xdc30 */
            {8'h00}, /* 0xdc2f */
            {8'h00}, /* 0xdc2e */
            {8'h00}, /* 0xdc2d */
            {8'h00}, /* 0xdc2c */
            {8'h00}, /* 0xdc2b */
            {8'h00}, /* 0xdc2a */
            {8'h00}, /* 0xdc29 */
            {8'h00}, /* 0xdc28 */
            {8'h00}, /* 0xdc27 */
            {8'h00}, /* 0xdc26 */
            {8'h00}, /* 0xdc25 */
            {8'h00}, /* 0xdc24 */
            {8'h00}, /* 0xdc23 */
            {8'h00}, /* 0xdc22 */
            {8'h00}, /* 0xdc21 */
            {8'h00}, /* 0xdc20 */
            {8'h00}, /* 0xdc1f */
            {8'h00}, /* 0xdc1e */
            {8'h00}, /* 0xdc1d */
            {8'h00}, /* 0xdc1c */
            {8'h00}, /* 0xdc1b */
            {8'h00}, /* 0xdc1a */
            {8'h00}, /* 0xdc19 */
            {8'h00}, /* 0xdc18 */
            {8'h00}, /* 0xdc17 */
            {8'h00}, /* 0xdc16 */
            {8'h00}, /* 0xdc15 */
            {8'h00}, /* 0xdc14 */
            {8'h00}, /* 0xdc13 */
            {8'h00}, /* 0xdc12 */
            {8'h00}, /* 0xdc11 */
            {8'h00}, /* 0xdc10 */
            {8'h00}, /* 0xdc0f */
            {8'h00}, /* 0xdc0e */
            {8'h00}, /* 0xdc0d */
            {8'h00}, /* 0xdc0c */
            {8'h00}, /* 0xdc0b */
            {8'h00}, /* 0xdc0a */
            {8'h00}, /* 0xdc09 */
            {8'h00}, /* 0xdc08 */
            {8'h00}, /* 0xdc07 */
            {8'h00}, /* 0xdc06 */
            {8'h00}, /* 0xdc05 */
            {8'h00}, /* 0xdc04 */
            {8'h00}, /* 0xdc03 */
            {8'h00}, /* 0xdc02 */
            {8'h00}, /* 0xdc01 */
            {8'h00}, /* 0xdc00 */
            {8'h00}, /* 0xdbff */
            {8'h00}, /* 0xdbfe */
            {8'h00}, /* 0xdbfd */
            {8'h00}, /* 0xdbfc */
            {8'h00}, /* 0xdbfb */
            {8'h00}, /* 0xdbfa */
            {8'h00}, /* 0xdbf9 */
            {8'h00}, /* 0xdbf8 */
            {8'h00}, /* 0xdbf7 */
            {8'h00}, /* 0xdbf6 */
            {8'h00}, /* 0xdbf5 */
            {8'h00}, /* 0xdbf4 */
            {8'h00}, /* 0xdbf3 */
            {8'h00}, /* 0xdbf2 */
            {8'h00}, /* 0xdbf1 */
            {8'h00}, /* 0xdbf0 */
            {8'h00}, /* 0xdbef */
            {8'h00}, /* 0xdbee */
            {8'h00}, /* 0xdbed */
            {8'h00}, /* 0xdbec */
            {8'h00}, /* 0xdbeb */
            {8'h00}, /* 0xdbea */
            {8'h00}, /* 0xdbe9 */
            {8'h00}, /* 0xdbe8 */
            {8'h00}, /* 0xdbe7 */
            {8'h00}, /* 0xdbe6 */
            {8'h00}, /* 0xdbe5 */
            {8'h00}, /* 0xdbe4 */
            {8'h00}, /* 0xdbe3 */
            {8'h00}, /* 0xdbe2 */
            {8'h00}, /* 0xdbe1 */
            {8'h00}, /* 0xdbe0 */
            {8'h00}, /* 0xdbdf */
            {8'h00}, /* 0xdbde */
            {8'h00}, /* 0xdbdd */
            {8'h00}, /* 0xdbdc */
            {8'h00}, /* 0xdbdb */
            {8'h00}, /* 0xdbda */
            {8'h00}, /* 0xdbd9 */
            {8'h00}, /* 0xdbd8 */
            {8'h00}, /* 0xdbd7 */
            {8'h00}, /* 0xdbd6 */
            {8'h00}, /* 0xdbd5 */
            {8'h00}, /* 0xdbd4 */
            {8'h00}, /* 0xdbd3 */
            {8'h00}, /* 0xdbd2 */
            {8'h00}, /* 0xdbd1 */
            {8'h00}, /* 0xdbd0 */
            {8'h00}, /* 0xdbcf */
            {8'h00}, /* 0xdbce */
            {8'h00}, /* 0xdbcd */
            {8'h00}, /* 0xdbcc */
            {8'h00}, /* 0xdbcb */
            {8'h00}, /* 0xdbca */
            {8'h00}, /* 0xdbc9 */
            {8'h00}, /* 0xdbc8 */
            {8'h00}, /* 0xdbc7 */
            {8'h00}, /* 0xdbc6 */
            {8'h00}, /* 0xdbc5 */
            {8'h00}, /* 0xdbc4 */
            {8'h00}, /* 0xdbc3 */
            {8'h00}, /* 0xdbc2 */
            {8'h00}, /* 0xdbc1 */
            {8'h00}, /* 0xdbc0 */
            {8'h00}, /* 0xdbbf */
            {8'h00}, /* 0xdbbe */
            {8'h00}, /* 0xdbbd */
            {8'h00}, /* 0xdbbc */
            {8'h00}, /* 0xdbbb */
            {8'h00}, /* 0xdbba */
            {8'h00}, /* 0xdbb9 */
            {8'h00}, /* 0xdbb8 */
            {8'h00}, /* 0xdbb7 */
            {8'h00}, /* 0xdbb6 */
            {8'h00}, /* 0xdbb5 */
            {8'h00}, /* 0xdbb4 */
            {8'h00}, /* 0xdbb3 */
            {8'h00}, /* 0xdbb2 */
            {8'h00}, /* 0xdbb1 */
            {8'h00}, /* 0xdbb0 */
            {8'h00}, /* 0xdbaf */
            {8'h00}, /* 0xdbae */
            {8'h00}, /* 0xdbad */
            {8'h00}, /* 0xdbac */
            {8'h00}, /* 0xdbab */
            {8'h00}, /* 0xdbaa */
            {8'h00}, /* 0xdba9 */
            {8'h00}, /* 0xdba8 */
            {8'h00}, /* 0xdba7 */
            {8'h00}, /* 0xdba6 */
            {8'h00}, /* 0xdba5 */
            {8'h00}, /* 0xdba4 */
            {8'h00}, /* 0xdba3 */
            {8'h00}, /* 0xdba2 */
            {8'h00}, /* 0xdba1 */
            {8'h00}, /* 0xdba0 */
            {8'h00}, /* 0xdb9f */
            {8'h00}, /* 0xdb9e */
            {8'h00}, /* 0xdb9d */
            {8'h00}, /* 0xdb9c */
            {8'h00}, /* 0xdb9b */
            {8'h00}, /* 0xdb9a */
            {8'h00}, /* 0xdb99 */
            {8'h00}, /* 0xdb98 */
            {8'h00}, /* 0xdb97 */
            {8'h00}, /* 0xdb96 */
            {8'h00}, /* 0xdb95 */
            {8'h00}, /* 0xdb94 */
            {8'h00}, /* 0xdb93 */
            {8'h00}, /* 0xdb92 */
            {8'h00}, /* 0xdb91 */
            {8'h00}, /* 0xdb90 */
            {8'h00}, /* 0xdb8f */
            {8'h00}, /* 0xdb8e */
            {8'h00}, /* 0xdb8d */
            {8'h00}, /* 0xdb8c */
            {8'h00}, /* 0xdb8b */
            {8'h00}, /* 0xdb8a */
            {8'h00}, /* 0xdb89 */
            {8'h00}, /* 0xdb88 */
            {8'h00}, /* 0xdb87 */
            {8'h00}, /* 0xdb86 */
            {8'h00}, /* 0xdb85 */
            {8'h00}, /* 0xdb84 */
            {8'h00}, /* 0xdb83 */
            {8'h00}, /* 0xdb82 */
            {8'h00}, /* 0xdb81 */
            {8'h00}, /* 0xdb80 */
            {8'h00}, /* 0xdb7f */
            {8'h00}, /* 0xdb7e */
            {8'h00}, /* 0xdb7d */
            {8'h00}, /* 0xdb7c */
            {8'h00}, /* 0xdb7b */
            {8'h00}, /* 0xdb7a */
            {8'h00}, /* 0xdb79 */
            {8'h00}, /* 0xdb78 */
            {8'h00}, /* 0xdb77 */
            {8'h00}, /* 0xdb76 */
            {8'h00}, /* 0xdb75 */
            {8'h00}, /* 0xdb74 */
            {8'h00}, /* 0xdb73 */
            {8'h00}, /* 0xdb72 */
            {8'h00}, /* 0xdb71 */
            {8'h00}, /* 0xdb70 */
            {8'h00}, /* 0xdb6f */
            {8'h00}, /* 0xdb6e */
            {8'h00}, /* 0xdb6d */
            {8'h00}, /* 0xdb6c */
            {8'h00}, /* 0xdb6b */
            {8'h00}, /* 0xdb6a */
            {8'h00}, /* 0xdb69 */
            {8'h00}, /* 0xdb68 */
            {8'h00}, /* 0xdb67 */
            {8'h00}, /* 0xdb66 */
            {8'h00}, /* 0xdb65 */
            {8'h00}, /* 0xdb64 */
            {8'h00}, /* 0xdb63 */
            {8'h00}, /* 0xdb62 */
            {8'h00}, /* 0xdb61 */
            {8'h00}, /* 0xdb60 */
            {8'h00}, /* 0xdb5f */
            {8'h00}, /* 0xdb5e */
            {8'h00}, /* 0xdb5d */
            {8'h00}, /* 0xdb5c */
            {8'h00}, /* 0xdb5b */
            {8'h00}, /* 0xdb5a */
            {8'h00}, /* 0xdb59 */
            {8'h00}, /* 0xdb58 */
            {8'h00}, /* 0xdb57 */
            {8'h00}, /* 0xdb56 */
            {8'h00}, /* 0xdb55 */
            {8'h00}, /* 0xdb54 */
            {8'h00}, /* 0xdb53 */
            {8'h00}, /* 0xdb52 */
            {8'h00}, /* 0xdb51 */
            {8'h00}, /* 0xdb50 */
            {8'h00}, /* 0xdb4f */
            {8'h00}, /* 0xdb4e */
            {8'h00}, /* 0xdb4d */
            {8'h00}, /* 0xdb4c */
            {8'h00}, /* 0xdb4b */
            {8'h00}, /* 0xdb4a */
            {8'h00}, /* 0xdb49 */
            {8'h00}, /* 0xdb48 */
            {8'h00}, /* 0xdb47 */
            {8'h00}, /* 0xdb46 */
            {8'h00}, /* 0xdb45 */
            {8'h00}, /* 0xdb44 */
            {8'h00}, /* 0xdb43 */
            {8'h00}, /* 0xdb42 */
            {8'h00}, /* 0xdb41 */
            {8'h00}, /* 0xdb40 */
            {8'h00}, /* 0xdb3f */
            {8'h00}, /* 0xdb3e */
            {8'h00}, /* 0xdb3d */
            {8'h00}, /* 0xdb3c */
            {8'h00}, /* 0xdb3b */
            {8'h00}, /* 0xdb3a */
            {8'h00}, /* 0xdb39 */
            {8'h00}, /* 0xdb38 */
            {8'h00}, /* 0xdb37 */
            {8'h00}, /* 0xdb36 */
            {8'h00}, /* 0xdb35 */
            {8'h00}, /* 0xdb34 */
            {8'h00}, /* 0xdb33 */
            {8'h00}, /* 0xdb32 */
            {8'h00}, /* 0xdb31 */
            {8'h00}, /* 0xdb30 */
            {8'h00}, /* 0xdb2f */
            {8'h00}, /* 0xdb2e */
            {8'h00}, /* 0xdb2d */
            {8'h00}, /* 0xdb2c */
            {8'h00}, /* 0xdb2b */
            {8'h00}, /* 0xdb2a */
            {8'h00}, /* 0xdb29 */
            {8'h00}, /* 0xdb28 */
            {8'h00}, /* 0xdb27 */
            {8'h00}, /* 0xdb26 */
            {8'h00}, /* 0xdb25 */
            {8'h00}, /* 0xdb24 */
            {8'h00}, /* 0xdb23 */
            {8'h00}, /* 0xdb22 */
            {8'h00}, /* 0xdb21 */
            {8'h00}, /* 0xdb20 */
            {8'h00}, /* 0xdb1f */
            {8'h00}, /* 0xdb1e */
            {8'h00}, /* 0xdb1d */
            {8'h00}, /* 0xdb1c */
            {8'h00}, /* 0xdb1b */
            {8'h00}, /* 0xdb1a */
            {8'h00}, /* 0xdb19 */
            {8'h00}, /* 0xdb18 */
            {8'h00}, /* 0xdb17 */
            {8'h00}, /* 0xdb16 */
            {8'h00}, /* 0xdb15 */
            {8'h00}, /* 0xdb14 */
            {8'h00}, /* 0xdb13 */
            {8'h00}, /* 0xdb12 */
            {8'h00}, /* 0xdb11 */
            {8'h00}, /* 0xdb10 */
            {8'h00}, /* 0xdb0f */
            {8'h00}, /* 0xdb0e */
            {8'h00}, /* 0xdb0d */
            {8'h00}, /* 0xdb0c */
            {8'h00}, /* 0xdb0b */
            {8'h00}, /* 0xdb0a */
            {8'h00}, /* 0xdb09 */
            {8'h00}, /* 0xdb08 */
            {8'h00}, /* 0xdb07 */
            {8'h00}, /* 0xdb06 */
            {8'h00}, /* 0xdb05 */
            {8'h00}, /* 0xdb04 */
            {8'h00}, /* 0xdb03 */
            {8'h00}, /* 0xdb02 */
            {8'h00}, /* 0xdb01 */
            {8'h00}, /* 0xdb00 */
            {8'h00}, /* 0xdaff */
            {8'h00}, /* 0xdafe */
            {8'h00}, /* 0xdafd */
            {8'h00}, /* 0xdafc */
            {8'h00}, /* 0xdafb */
            {8'h00}, /* 0xdafa */
            {8'h00}, /* 0xdaf9 */
            {8'h00}, /* 0xdaf8 */
            {8'h00}, /* 0xdaf7 */
            {8'h00}, /* 0xdaf6 */
            {8'h00}, /* 0xdaf5 */
            {8'h00}, /* 0xdaf4 */
            {8'h00}, /* 0xdaf3 */
            {8'h00}, /* 0xdaf2 */
            {8'h00}, /* 0xdaf1 */
            {8'h00}, /* 0xdaf0 */
            {8'h00}, /* 0xdaef */
            {8'h00}, /* 0xdaee */
            {8'h00}, /* 0xdaed */
            {8'h00}, /* 0xdaec */
            {8'h00}, /* 0xdaeb */
            {8'h00}, /* 0xdaea */
            {8'h00}, /* 0xdae9 */
            {8'h00}, /* 0xdae8 */
            {8'h00}, /* 0xdae7 */
            {8'h00}, /* 0xdae6 */
            {8'h00}, /* 0xdae5 */
            {8'h00}, /* 0xdae4 */
            {8'h00}, /* 0xdae3 */
            {8'h00}, /* 0xdae2 */
            {8'h00}, /* 0xdae1 */
            {8'h00}, /* 0xdae0 */
            {8'h00}, /* 0xdadf */
            {8'h00}, /* 0xdade */
            {8'h00}, /* 0xdadd */
            {8'h00}, /* 0xdadc */
            {8'h00}, /* 0xdadb */
            {8'h00}, /* 0xdada */
            {8'h00}, /* 0xdad9 */
            {8'h00}, /* 0xdad8 */
            {8'h00}, /* 0xdad7 */
            {8'h00}, /* 0xdad6 */
            {8'h00}, /* 0xdad5 */
            {8'h00}, /* 0xdad4 */
            {8'h00}, /* 0xdad3 */
            {8'h00}, /* 0xdad2 */
            {8'h00}, /* 0xdad1 */
            {8'h00}, /* 0xdad0 */
            {8'h00}, /* 0xdacf */
            {8'h00}, /* 0xdace */
            {8'h00}, /* 0xdacd */
            {8'h00}, /* 0xdacc */
            {8'h00}, /* 0xdacb */
            {8'h00}, /* 0xdaca */
            {8'h00}, /* 0xdac9 */
            {8'h00}, /* 0xdac8 */
            {8'h00}, /* 0xdac7 */
            {8'h00}, /* 0xdac6 */
            {8'h00}, /* 0xdac5 */
            {8'h00}, /* 0xdac4 */
            {8'h00}, /* 0xdac3 */
            {8'h00}, /* 0xdac2 */
            {8'h00}, /* 0xdac1 */
            {8'h00}, /* 0xdac0 */
            {8'h00}, /* 0xdabf */
            {8'h00}, /* 0xdabe */
            {8'h00}, /* 0xdabd */
            {8'h00}, /* 0xdabc */
            {8'h00}, /* 0xdabb */
            {8'h00}, /* 0xdaba */
            {8'h00}, /* 0xdab9 */
            {8'h00}, /* 0xdab8 */
            {8'h00}, /* 0xdab7 */
            {8'h00}, /* 0xdab6 */
            {8'h00}, /* 0xdab5 */
            {8'h00}, /* 0xdab4 */
            {8'h00}, /* 0xdab3 */
            {8'h00}, /* 0xdab2 */
            {8'h00}, /* 0xdab1 */
            {8'h00}, /* 0xdab0 */
            {8'h00}, /* 0xdaaf */
            {8'h00}, /* 0xdaae */
            {8'h00}, /* 0xdaad */
            {8'h00}, /* 0xdaac */
            {8'h00}, /* 0xdaab */
            {8'h00}, /* 0xdaaa */
            {8'h00}, /* 0xdaa9 */
            {8'h00}, /* 0xdaa8 */
            {8'h00}, /* 0xdaa7 */
            {8'h00}, /* 0xdaa6 */
            {8'h00}, /* 0xdaa5 */
            {8'h00}, /* 0xdaa4 */
            {8'h00}, /* 0xdaa3 */
            {8'h00}, /* 0xdaa2 */
            {8'h00}, /* 0xdaa1 */
            {8'h00}, /* 0xdaa0 */
            {8'h00}, /* 0xda9f */
            {8'h00}, /* 0xda9e */
            {8'h00}, /* 0xda9d */
            {8'h00}, /* 0xda9c */
            {8'h00}, /* 0xda9b */
            {8'h00}, /* 0xda9a */
            {8'h00}, /* 0xda99 */
            {8'h00}, /* 0xda98 */
            {8'h00}, /* 0xda97 */
            {8'h00}, /* 0xda96 */
            {8'h00}, /* 0xda95 */
            {8'h00}, /* 0xda94 */
            {8'h00}, /* 0xda93 */
            {8'h00}, /* 0xda92 */
            {8'h00}, /* 0xda91 */
            {8'h00}, /* 0xda90 */
            {8'h00}, /* 0xda8f */
            {8'h00}, /* 0xda8e */
            {8'h00}, /* 0xda8d */
            {8'h00}, /* 0xda8c */
            {8'h00}, /* 0xda8b */
            {8'h00}, /* 0xda8a */
            {8'h00}, /* 0xda89 */
            {8'h00}, /* 0xda88 */
            {8'h00}, /* 0xda87 */
            {8'h00}, /* 0xda86 */
            {8'h00}, /* 0xda85 */
            {8'h00}, /* 0xda84 */
            {8'h00}, /* 0xda83 */
            {8'h00}, /* 0xda82 */
            {8'h00}, /* 0xda81 */
            {8'h00}, /* 0xda80 */
            {8'h00}, /* 0xda7f */
            {8'h00}, /* 0xda7e */
            {8'h00}, /* 0xda7d */
            {8'h00}, /* 0xda7c */
            {8'h00}, /* 0xda7b */
            {8'h00}, /* 0xda7a */
            {8'h00}, /* 0xda79 */
            {8'h00}, /* 0xda78 */
            {8'h00}, /* 0xda77 */
            {8'h00}, /* 0xda76 */
            {8'h00}, /* 0xda75 */
            {8'h00}, /* 0xda74 */
            {8'h00}, /* 0xda73 */
            {8'h00}, /* 0xda72 */
            {8'h00}, /* 0xda71 */
            {8'h00}, /* 0xda70 */
            {8'h00}, /* 0xda6f */
            {8'h00}, /* 0xda6e */
            {8'h00}, /* 0xda6d */
            {8'h00}, /* 0xda6c */
            {8'h00}, /* 0xda6b */
            {8'h00}, /* 0xda6a */
            {8'h00}, /* 0xda69 */
            {8'h00}, /* 0xda68 */
            {8'h00}, /* 0xda67 */
            {8'h00}, /* 0xda66 */
            {8'h00}, /* 0xda65 */
            {8'h00}, /* 0xda64 */
            {8'h00}, /* 0xda63 */
            {8'h00}, /* 0xda62 */
            {8'h00}, /* 0xda61 */
            {8'h00}, /* 0xda60 */
            {8'h00}, /* 0xda5f */
            {8'h00}, /* 0xda5e */
            {8'h00}, /* 0xda5d */
            {8'h00}, /* 0xda5c */
            {8'h00}, /* 0xda5b */
            {8'h00}, /* 0xda5a */
            {8'h00}, /* 0xda59 */
            {8'h00}, /* 0xda58 */
            {8'h00}, /* 0xda57 */
            {8'h00}, /* 0xda56 */
            {8'h00}, /* 0xda55 */
            {8'h00}, /* 0xda54 */
            {8'h00}, /* 0xda53 */
            {8'h00}, /* 0xda52 */
            {8'h00}, /* 0xda51 */
            {8'h00}, /* 0xda50 */
            {8'h00}, /* 0xda4f */
            {8'h00}, /* 0xda4e */
            {8'h00}, /* 0xda4d */
            {8'h00}, /* 0xda4c */
            {8'h00}, /* 0xda4b */
            {8'h00}, /* 0xda4a */
            {8'h00}, /* 0xda49 */
            {8'h00}, /* 0xda48 */
            {8'h00}, /* 0xda47 */
            {8'h00}, /* 0xda46 */
            {8'h00}, /* 0xda45 */
            {8'h00}, /* 0xda44 */
            {8'h00}, /* 0xda43 */
            {8'h00}, /* 0xda42 */
            {8'h00}, /* 0xda41 */
            {8'h00}, /* 0xda40 */
            {8'h00}, /* 0xda3f */
            {8'h00}, /* 0xda3e */
            {8'h00}, /* 0xda3d */
            {8'h00}, /* 0xda3c */
            {8'h00}, /* 0xda3b */
            {8'h00}, /* 0xda3a */
            {8'h00}, /* 0xda39 */
            {8'h00}, /* 0xda38 */
            {8'h00}, /* 0xda37 */
            {8'h00}, /* 0xda36 */
            {8'h00}, /* 0xda35 */
            {8'h00}, /* 0xda34 */
            {8'h00}, /* 0xda33 */
            {8'h00}, /* 0xda32 */
            {8'h00}, /* 0xda31 */
            {8'h00}, /* 0xda30 */
            {8'h00}, /* 0xda2f */
            {8'h00}, /* 0xda2e */
            {8'h00}, /* 0xda2d */
            {8'h00}, /* 0xda2c */
            {8'h00}, /* 0xda2b */
            {8'h00}, /* 0xda2a */
            {8'h00}, /* 0xda29 */
            {8'h00}, /* 0xda28 */
            {8'h00}, /* 0xda27 */
            {8'h00}, /* 0xda26 */
            {8'h00}, /* 0xda25 */
            {8'h00}, /* 0xda24 */
            {8'h00}, /* 0xda23 */
            {8'h00}, /* 0xda22 */
            {8'h00}, /* 0xda21 */
            {8'h00}, /* 0xda20 */
            {8'h00}, /* 0xda1f */
            {8'h00}, /* 0xda1e */
            {8'h00}, /* 0xda1d */
            {8'h00}, /* 0xda1c */
            {8'h00}, /* 0xda1b */
            {8'h00}, /* 0xda1a */
            {8'h00}, /* 0xda19 */
            {8'h00}, /* 0xda18 */
            {8'h00}, /* 0xda17 */
            {8'h00}, /* 0xda16 */
            {8'h00}, /* 0xda15 */
            {8'h00}, /* 0xda14 */
            {8'h00}, /* 0xda13 */
            {8'h00}, /* 0xda12 */
            {8'h00}, /* 0xda11 */
            {8'h00}, /* 0xda10 */
            {8'h00}, /* 0xda0f */
            {8'h00}, /* 0xda0e */
            {8'h00}, /* 0xda0d */
            {8'h00}, /* 0xda0c */
            {8'h00}, /* 0xda0b */
            {8'h00}, /* 0xda0a */
            {8'h00}, /* 0xda09 */
            {8'h00}, /* 0xda08 */
            {8'h00}, /* 0xda07 */
            {8'h00}, /* 0xda06 */
            {8'h00}, /* 0xda05 */
            {8'h00}, /* 0xda04 */
            {8'h00}, /* 0xda03 */
            {8'h00}, /* 0xda02 */
            {8'h00}, /* 0xda01 */
            {8'h00}, /* 0xda00 */
            {8'h00}, /* 0xd9ff */
            {8'h00}, /* 0xd9fe */
            {8'h00}, /* 0xd9fd */
            {8'h00}, /* 0xd9fc */
            {8'h00}, /* 0xd9fb */
            {8'h00}, /* 0xd9fa */
            {8'h00}, /* 0xd9f9 */
            {8'h00}, /* 0xd9f8 */
            {8'h00}, /* 0xd9f7 */
            {8'h00}, /* 0xd9f6 */
            {8'h00}, /* 0xd9f5 */
            {8'h00}, /* 0xd9f4 */
            {8'h00}, /* 0xd9f3 */
            {8'h00}, /* 0xd9f2 */
            {8'h00}, /* 0xd9f1 */
            {8'h00}, /* 0xd9f0 */
            {8'h00}, /* 0xd9ef */
            {8'h00}, /* 0xd9ee */
            {8'h00}, /* 0xd9ed */
            {8'h00}, /* 0xd9ec */
            {8'h00}, /* 0xd9eb */
            {8'h00}, /* 0xd9ea */
            {8'h00}, /* 0xd9e9 */
            {8'h00}, /* 0xd9e8 */
            {8'h00}, /* 0xd9e7 */
            {8'h00}, /* 0xd9e6 */
            {8'h00}, /* 0xd9e5 */
            {8'h00}, /* 0xd9e4 */
            {8'h00}, /* 0xd9e3 */
            {8'h00}, /* 0xd9e2 */
            {8'h00}, /* 0xd9e1 */
            {8'h00}, /* 0xd9e0 */
            {8'h00}, /* 0xd9df */
            {8'h00}, /* 0xd9de */
            {8'h00}, /* 0xd9dd */
            {8'h00}, /* 0xd9dc */
            {8'h00}, /* 0xd9db */
            {8'h00}, /* 0xd9da */
            {8'h00}, /* 0xd9d9 */
            {8'h00}, /* 0xd9d8 */
            {8'h00}, /* 0xd9d7 */
            {8'h00}, /* 0xd9d6 */
            {8'h00}, /* 0xd9d5 */
            {8'h00}, /* 0xd9d4 */
            {8'h00}, /* 0xd9d3 */
            {8'h00}, /* 0xd9d2 */
            {8'h00}, /* 0xd9d1 */
            {8'h00}, /* 0xd9d0 */
            {8'h00}, /* 0xd9cf */
            {8'h00}, /* 0xd9ce */
            {8'h00}, /* 0xd9cd */
            {8'h00}, /* 0xd9cc */
            {8'h00}, /* 0xd9cb */
            {8'h00}, /* 0xd9ca */
            {8'h00}, /* 0xd9c9 */
            {8'h00}, /* 0xd9c8 */
            {8'h00}, /* 0xd9c7 */
            {8'h00}, /* 0xd9c6 */
            {8'h00}, /* 0xd9c5 */
            {8'h00}, /* 0xd9c4 */
            {8'h00}, /* 0xd9c3 */
            {8'h00}, /* 0xd9c2 */
            {8'h00}, /* 0xd9c1 */
            {8'h00}, /* 0xd9c0 */
            {8'h00}, /* 0xd9bf */
            {8'h00}, /* 0xd9be */
            {8'h00}, /* 0xd9bd */
            {8'h00}, /* 0xd9bc */
            {8'h00}, /* 0xd9bb */
            {8'h00}, /* 0xd9ba */
            {8'h00}, /* 0xd9b9 */
            {8'h00}, /* 0xd9b8 */
            {8'h00}, /* 0xd9b7 */
            {8'h00}, /* 0xd9b6 */
            {8'h00}, /* 0xd9b5 */
            {8'h00}, /* 0xd9b4 */
            {8'h00}, /* 0xd9b3 */
            {8'h00}, /* 0xd9b2 */
            {8'h00}, /* 0xd9b1 */
            {8'h00}, /* 0xd9b0 */
            {8'h00}, /* 0xd9af */
            {8'h00}, /* 0xd9ae */
            {8'h00}, /* 0xd9ad */
            {8'h00}, /* 0xd9ac */
            {8'h00}, /* 0xd9ab */
            {8'h00}, /* 0xd9aa */
            {8'h00}, /* 0xd9a9 */
            {8'h00}, /* 0xd9a8 */
            {8'h00}, /* 0xd9a7 */
            {8'h00}, /* 0xd9a6 */
            {8'h00}, /* 0xd9a5 */
            {8'h00}, /* 0xd9a4 */
            {8'h00}, /* 0xd9a3 */
            {8'h00}, /* 0xd9a2 */
            {8'h00}, /* 0xd9a1 */
            {8'h00}, /* 0xd9a0 */
            {8'h00}, /* 0xd99f */
            {8'h00}, /* 0xd99e */
            {8'h00}, /* 0xd99d */
            {8'h00}, /* 0xd99c */
            {8'h00}, /* 0xd99b */
            {8'h00}, /* 0xd99a */
            {8'h00}, /* 0xd999 */
            {8'h00}, /* 0xd998 */
            {8'h00}, /* 0xd997 */
            {8'h00}, /* 0xd996 */
            {8'h00}, /* 0xd995 */
            {8'h00}, /* 0xd994 */
            {8'h00}, /* 0xd993 */
            {8'h00}, /* 0xd992 */
            {8'h00}, /* 0xd991 */
            {8'h00}, /* 0xd990 */
            {8'h00}, /* 0xd98f */
            {8'h00}, /* 0xd98e */
            {8'h00}, /* 0xd98d */
            {8'h00}, /* 0xd98c */
            {8'h00}, /* 0xd98b */
            {8'h00}, /* 0xd98a */
            {8'h00}, /* 0xd989 */
            {8'h00}, /* 0xd988 */
            {8'h00}, /* 0xd987 */
            {8'h00}, /* 0xd986 */
            {8'h00}, /* 0xd985 */
            {8'h00}, /* 0xd984 */
            {8'h00}, /* 0xd983 */
            {8'h00}, /* 0xd982 */
            {8'h00}, /* 0xd981 */
            {8'h00}, /* 0xd980 */
            {8'h00}, /* 0xd97f */
            {8'h00}, /* 0xd97e */
            {8'h00}, /* 0xd97d */
            {8'h00}, /* 0xd97c */
            {8'h00}, /* 0xd97b */
            {8'h00}, /* 0xd97a */
            {8'h00}, /* 0xd979 */
            {8'h00}, /* 0xd978 */
            {8'h00}, /* 0xd977 */
            {8'h00}, /* 0xd976 */
            {8'h00}, /* 0xd975 */
            {8'h00}, /* 0xd974 */
            {8'h00}, /* 0xd973 */
            {8'h00}, /* 0xd972 */
            {8'h00}, /* 0xd971 */
            {8'h00}, /* 0xd970 */
            {8'h00}, /* 0xd96f */
            {8'h00}, /* 0xd96e */
            {8'h00}, /* 0xd96d */
            {8'h00}, /* 0xd96c */
            {8'h00}, /* 0xd96b */
            {8'h00}, /* 0xd96a */
            {8'h00}, /* 0xd969 */
            {8'h00}, /* 0xd968 */
            {8'h00}, /* 0xd967 */
            {8'h00}, /* 0xd966 */
            {8'h00}, /* 0xd965 */
            {8'h00}, /* 0xd964 */
            {8'h00}, /* 0xd963 */
            {8'h00}, /* 0xd962 */
            {8'h00}, /* 0xd961 */
            {8'h00}, /* 0xd960 */
            {8'h00}, /* 0xd95f */
            {8'h00}, /* 0xd95e */
            {8'h00}, /* 0xd95d */
            {8'h00}, /* 0xd95c */
            {8'h00}, /* 0xd95b */
            {8'h00}, /* 0xd95a */
            {8'h00}, /* 0xd959 */
            {8'h00}, /* 0xd958 */
            {8'h00}, /* 0xd957 */
            {8'h00}, /* 0xd956 */
            {8'h00}, /* 0xd955 */
            {8'h00}, /* 0xd954 */
            {8'h00}, /* 0xd953 */
            {8'h00}, /* 0xd952 */
            {8'h00}, /* 0xd951 */
            {8'h00}, /* 0xd950 */
            {8'h00}, /* 0xd94f */
            {8'h00}, /* 0xd94e */
            {8'h00}, /* 0xd94d */
            {8'h00}, /* 0xd94c */
            {8'h00}, /* 0xd94b */
            {8'h00}, /* 0xd94a */
            {8'h00}, /* 0xd949 */
            {8'h00}, /* 0xd948 */
            {8'h00}, /* 0xd947 */
            {8'h00}, /* 0xd946 */
            {8'h00}, /* 0xd945 */
            {8'h00}, /* 0xd944 */
            {8'h00}, /* 0xd943 */
            {8'h00}, /* 0xd942 */
            {8'h00}, /* 0xd941 */
            {8'h00}, /* 0xd940 */
            {8'h00}, /* 0xd93f */
            {8'h00}, /* 0xd93e */
            {8'h00}, /* 0xd93d */
            {8'h00}, /* 0xd93c */
            {8'h00}, /* 0xd93b */
            {8'h00}, /* 0xd93a */
            {8'h00}, /* 0xd939 */
            {8'h00}, /* 0xd938 */
            {8'h00}, /* 0xd937 */
            {8'h00}, /* 0xd936 */
            {8'h00}, /* 0xd935 */
            {8'h00}, /* 0xd934 */
            {8'h00}, /* 0xd933 */
            {8'h00}, /* 0xd932 */
            {8'h00}, /* 0xd931 */
            {8'h00}, /* 0xd930 */
            {8'h00}, /* 0xd92f */
            {8'h00}, /* 0xd92e */
            {8'h00}, /* 0xd92d */
            {8'h00}, /* 0xd92c */
            {8'h00}, /* 0xd92b */
            {8'h00}, /* 0xd92a */
            {8'h00}, /* 0xd929 */
            {8'h00}, /* 0xd928 */
            {8'h00}, /* 0xd927 */
            {8'h00}, /* 0xd926 */
            {8'h00}, /* 0xd925 */
            {8'h00}, /* 0xd924 */
            {8'h00}, /* 0xd923 */
            {8'h00}, /* 0xd922 */
            {8'h00}, /* 0xd921 */
            {8'h00}, /* 0xd920 */
            {8'h00}, /* 0xd91f */
            {8'h00}, /* 0xd91e */
            {8'h00}, /* 0xd91d */
            {8'h00}, /* 0xd91c */
            {8'h00}, /* 0xd91b */
            {8'h00}, /* 0xd91a */
            {8'h00}, /* 0xd919 */
            {8'h00}, /* 0xd918 */
            {8'h00}, /* 0xd917 */
            {8'h00}, /* 0xd916 */
            {8'h00}, /* 0xd915 */
            {8'h00}, /* 0xd914 */
            {8'h00}, /* 0xd913 */
            {8'h00}, /* 0xd912 */
            {8'h00}, /* 0xd911 */
            {8'h00}, /* 0xd910 */
            {8'h00}, /* 0xd90f */
            {8'h00}, /* 0xd90e */
            {8'h00}, /* 0xd90d */
            {8'h00}, /* 0xd90c */
            {8'h00}, /* 0xd90b */
            {8'h00}, /* 0xd90a */
            {8'h00}, /* 0xd909 */
            {8'h00}, /* 0xd908 */
            {8'h00}, /* 0xd907 */
            {8'h00}, /* 0xd906 */
            {8'h00}, /* 0xd905 */
            {8'h00}, /* 0xd904 */
            {8'h00}, /* 0xd903 */
            {8'h00}, /* 0xd902 */
            {8'h00}, /* 0xd901 */
            {8'h00}, /* 0xd900 */
            {8'h00}, /* 0xd8ff */
            {8'h00}, /* 0xd8fe */
            {8'h00}, /* 0xd8fd */
            {8'h00}, /* 0xd8fc */
            {8'h00}, /* 0xd8fb */
            {8'h00}, /* 0xd8fa */
            {8'h00}, /* 0xd8f9 */
            {8'h00}, /* 0xd8f8 */
            {8'h00}, /* 0xd8f7 */
            {8'h00}, /* 0xd8f6 */
            {8'h00}, /* 0xd8f5 */
            {8'h00}, /* 0xd8f4 */
            {8'h00}, /* 0xd8f3 */
            {8'h00}, /* 0xd8f2 */
            {8'h00}, /* 0xd8f1 */
            {8'h00}, /* 0xd8f0 */
            {8'h00}, /* 0xd8ef */
            {8'h00}, /* 0xd8ee */
            {8'h00}, /* 0xd8ed */
            {8'h00}, /* 0xd8ec */
            {8'h00}, /* 0xd8eb */
            {8'h00}, /* 0xd8ea */
            {8'h00}, /* 0xd8e9 */
            {8'h00}, /* 0xd8e8 */
            {8'h00}, /* 0xd8e7 */
            {8'h00}, /* 0xd8e6 */
            {8'h00}, /* 0xd8e5 */
            {8'h00}, /* 0xd8e4 */
            {8'h00}, /* 0xd8e3 */
            {8'h00}, /* 0xd8e2 */
            {8'h00}, /* 0xd8e1 */
            {8'h00}, /* 0xd8e0 */
            {8'h00}, /* 0xd8df */
            {8'h00}, /* 0xd8de */
            {8'h00}, /* 0xd8dd */
            {8'h00}, /* 0xd8dc */
            {8'h00}, /* 0xd8db */
            {8'h00}, /* 0xd8da */
            {8'h00}, /* 0xd8d9 */
            {8'h00}, /* 0xd8d8 */
            {8'h00}, /* 0xd8d7 */
            {8'h00}, /* 0xd8d6 */
            {8'h00}, /* 0xd8d5 */
            {8'h00}, /* 0xd8d4 */
            {8'h00}, /* 0xd8d3 */
            {8'h00}, /* 0xd8d2 */
            {8'h00}, /* 0xd8d1 */
            {8'h00}, /* 0xd8d0 */
            {8'h00}, /* 0xd8cf */
            {8'h00}, /* 0xd8ce */
            {8'h00}, /* 0xd8cd */
            {8'h00}, /* 0xd8cc */
            {8'h00}, /* 0xd8cb */
            {8'h00}, /* 0xd8ca */
            {8'h00}, /* 0xd8c9 */
            {8'h00}, /* 0xd8c8 */
            {8'h00}, /* 0xd8c7 */
            {8'h00}, /* 0xd8c6 */
            {8'h00}, /* 0xd8c5 */
            {8'h00}, /* 0xd8c4 */
            {8'h00}, /* 0xd8c3 */
            {8'h00}, /* 0xd8c2 */
            {8'h00}, /* 0xd8c1 */
            {8'h00}, /* 0xd8c0 */
            {8'h00}, /* 0xd8bf */
            {8'h00}, /* 0xd8be */
            {8'h00}, /* 0xd8bd */
            {8'h00}, /* 0xd8bc */
            {8'h00}, /* 0xd8bb */
            {8'h00}, /* 0xd8ba */
            {8'h00}, /* 0xd8b9 */
            {8'h00}, /* 0xd8b8 */
            {8'h00}, /* 0xd8b7 */
            {8'h00}, /* 0xd8b6 */
            {8'h00}, /* 0xd8b5 */
            {8'h00}, /* 0xd8b4 */
            {8'h00}, /* 0xd8b3 */
            {8'h00}, /* 0xd8b2 */
            {8'h00}, /* 0xd8b1 */
            {8'h00}, /* 0xd8b0 */
            {8'h00}, /* 0xd8af */
            {8'h00}, /* 0xd8ae */
            {8'h00}, /* 0xd8ad */
            {8'h00}, /* 0xd8ac */
            {8'h00}, /* 0xd8ab */
            {8'h00}, /* 0xd8aa */
            {8'h00}, /* 0xd8a9 */
            {8'h00}, /* 0xd8a8 */
            {8'h00}, /* 0xd8a7 */
            {8'h00}, /* 0xd8a6 */
            {8'h00}, /* 0xd8a5 */
            {8'h00}, /* 0xd8a4 */
            {8'h00}, /* 0xd8a3 */
            {8'h00}, /* 0xd8a2 */
            {8'h00}, /* 0xd8a1 */
            {8'h00}, /* 0xd8a0 */
            {8'h00}, /* 0xd89f */
            {8'h00}, /* 0xd89e */
            {8'h00}, /* 0xd89d */
            {8'h00}, /* 0xd89c */
            {8'h00}, /* 0xd89b */
            {8'h00}, /* 0xd89a */
            {8'h00}, /* 0xd899 */
            {8'h00}, /* 0xd898 */
            {8'h00}, /* 0xd897 */
            {8'h00}, /* 0xd896 */
            {8'h00}, /* 0xd895 */
            {8'h00}, /* 0xd894 */
            {8'h00}, /* 0xd893 */
            {8'h00}, /* 0xd892 */
            {8'h00}, /* 0xd891 */
            {8'h00}, /* 0xd890 */
            {8'h00}, /* 0xd88f */
            {8'h00}, /* 0xd88e */
            {8'h00}, /* 0xd88d */
            {8'h00}, /* 0xd88c */
            {8'h00}, /* 0xd88b */
            {8'h00}, /* 0xd88a */
            {8'h00}, /* 0xd889 */
            {8'h00}, /* 0xd888 */
            {8'h00}, /* 0xd887 */
            {8'h00}, /* 0xd886 */
            {8'h00}, /* 0xd885 */
            {8'h00}, /* 0xd884 */
            {8'h00}, /* 0xd883 */
            {8'h00}, /* 0xd882 */
            {8'h00}, /* 0xd881 */
            {8'h00}, /* 0xd880 */
            {8'h00}, /* 0xd87f */
            {8'h00}, /* 0xd87e */
            {8'h00}, /* 0xd87d */
            {8'h00}, /* 0xd87c */
            {8'h00}, /* 0xd87b */
            {8'h00}, /* 0xd87a */
            {8'h00}, /* 0xd879 */
            {8'h00}, /* 0xd878 */
            {8'h00}, /* 0xd877 */
            {8'h00}, /* 0xd876 */
            {8'h00}, /* 0xd875 */
            {8'h00}, /* 0xd874 */
            {8'h00}, /* 0xd873 */
            {8'h00}, /* 0xd872 */
            {8'h00}, /* 0xd871 */
            {8'h00}, /* 0xd870 */
            {8'h00}, /* 0xd86f */
            {8'h00}, /* 0xd86e */
            {8'h00}, /* 0xd86d */
            {8'h00}, /* 0xd86c */
            {8'h00}, /* 0xd86b */
            {8'h00}, /* 0xd86a */
            {8'h00}, /* 0xd869 */
            {8'h00}, /* 0xd868 */
            {8'h00}, /* 0xd867 */
            {8'h00}, /* 0xd866 */
            {8'h00}, /* 0xd865 */
            {8'h00}, /* 0xd864 */
            {8'h00}, /* 0xd863 */
            {8'h00}, /* 0xd862 */
            {8'h00}, /* 0xd861 */
            {8'h00}, /* 0xd860 */
            {8'h00}, /* 0xd85f */
            {8'h00}, /* 0xd85e */
            {8'h00}, /* 0xd85d */
            {8'h00}, /* 0xd85c */
            {8'h00}, /* 0xd85b */
            {8'h00}, /* 0xd85a */
            {8'h00}, /* 0xd859 */
            {8'h00}, /* 0xd858 */
            {8'h00}, /* 0xd857 */
            {8'h00}, /* 0xd856 */
            {8'h00}, /* 0xd855 */
            {8'h00}, /* 0xd854 */
            {8'h00}, /* 0xd853 */
            {8'h00}, /* 0xd852 */
            {8'h00}, /* 0xd851 */
            {8'h00}, /* 0xd850 */
            {8'h00}, /* 0xd84f */
            {8'h00}, /* 0xd84e */
            {8'h00}, /* 0xd84d */
            {8'h00}, /* 0xd84c */
            {8'h00}, /* 0xd84b */
            {8'h00}, /* 0xd84a */
            {8'h00}, /* 0xd849 */
            {8'h00}, /* 0xd848 */
            {8'h00}, /* 0xd847 */
            {8'h00}, /* 0xd846 */
            {8'h00}, /* 0xd845 */
            {8'h00}, /* 0xd844 */
            {8'h00}, /* 0xd843 */
            {8'h00}, /* 0xd842 */
            {8'h00}, /* 0xd841 */
            {8'h00}, /* 0xd840 */
            {8'h00}, /* 0xd83f */
            {8'h00}, /* 0xd83e */
            {8'h00}, /* 0xd83d */
            {8'h00}, /* 0xd83c */
            {8'h00}, /* 0xd83b */
            {8'h00}, /* 0xd83a */
            {8'h00}, /* 0xd839 */
            {8'h00}, /* 0xd838 */
            {8'h00}, /* 0xd837 */
            {8'h00}, /* 0xd836 */
            {8'h00}, /* 0xd835 */
            {8'h00}, /* 0xd834 */
            {8'h00}, /* 0xd833 */
            {8'h00}, /* 0xd832 */
            {8'h00}, /* 0xd831 */
            {8'h00}, /* 0xd830 */
            {8'h00}, /* 0xd82f */
            {8'h00}, /* 0xd82e */
            {8'h00}, /* 0xd82d */
            {8'h00}, /* 0xd82c */
            {8'h00}, /* 0xd82b */
            {8'h00}, /* 0xd82a */
            {8'h00}, /* 0xd829 */
            {8'h00}, /* 0xd828 */
            {8'h00}, /* 0xd827 */
            {8'h00}, /* 0xd826 */
            {8'h00}, /* 0xd825 */
            {8'h00}, /* 0xd824 */
            {8'h00}, /* 0xd823 */
            {8'h00}, /* 0xd822 */
            {8'h00}, /* 0xd821 */
            {8'h00}, /* 0xd820 */
            {8'h00}, /* 0xd81f */
            {8'h00}, /* 0xd81e */
            {8'h00}, /* 0xd81d */
            {8'h00}, /* 0xd81c */
            {8'h00}, /* 0xd81b */
            {8'h00}, /* 0xd81a */
            {8'h00}, /* 0xd819 */
            {8'h00}, /* 0xd818 */
            {8'h00}, /* 0xd817 */
            {8'h00}, /* 0xd816 */
            {8'h00}, /* 0xd815 */
            {8'h00}, /* 0xd814 */
            {8'h00}, /* 0xd813 */
            {8'h00}, /* 0xd812 */
            {8'h00}, /* 0xd811 */
            {8'h00}, /* 0xd810 */
            {8'h00}, /* 0xd80f */
            {8'h00}, /* 0xd80e */
            {8'h00}, /* 0xd80d */
            {8'h00}, /* 0xd80c */
            {8'h00}, /* 0xd80b */
            {8'h00}, /* 0xd80a */
            {8'h00}, /* 0xd809 */
            {8'h00}, /* 0xd808 */
            {8'h00}, /* 0xd807 */
            {8'h00}, /* 0xd806 */
            {8'h00}, /* 0xd805 */
            {8'h00}, /* 0xd804 */
            {8'h00}, /* 0xd803 */
            {8'h00}, /* 0xd802 */
            {8'h00}, /* 0xd801 */
            {8'h00}, /* 0xd800 */
            {8'h00}, /* 0xd7ff */
            {8'h00}, /* 0xd7fe */
            {8'h00}, /* 0xd7fd */
            {8'h00}, /* 0xd7fc */
            {8'h00}, /* 0xd7fb */
            {8'h00}, /* 0xd7fa */
            {8'h00}, /* 0xd7f9 */
            {8'h00}, /* 0xd7f8 */
            {8'h00}, /* 0xd7f7 */
            {8'h00}, /* 0xd7f6 */
            {8'h00}, /* 0xd7f5 */
            {8'h00}, /* 0xd7f4 */
            {8'h00}, /* 0xd7f3 */
            {8'h00}, /* 0xd7f2 */
            {8'h00}, /* 0xd7f1 */
            {8'h00}, /* 0xd7f0 */
            {8'h00}, /* 0xd7ef */
            {8'h00}, /* 0xd7ee */
            {8'h00}, /* 0xd7ed */
            {8'h00}, /* 0xd7ec */
            {8'h00}, /* 0xd7eb */
            {8'h00}, /* 0xd7ea */
            {8'h00}, /* 0xd7e9 */
            {8'h00}, /* 0xd7e8 */
            {8'h00}, /* 0xd7e7 */
            {8'h00}, /* 0xd7e6 */
            {8'h00}, /* 0xd7e5 */
            {8'h00}, /* 0xd7e4 */
            {8'h00}, /* 0xd7e3 */
            {8'h00}, /* 0xd7e2 */
            {8'h00}, /* 0xd7e1 */
            {8'h00}, /* 0xd7e0 */
            {8'h00}, /* 0xd7df */
            {8'h00}, /* 0xd7de */
            {8'h00}, /* 0xd7dd */
            {8'h00}, /* 0xd7dc */
            {8'h00}, /* 0xd7db */
            {8'h00}, /* 0xd7da */
            {8'h00}, /* 0xd7d9 */
            {8'h00}, /* 0xd7d8 */
            {8'h00}, /* 0xd7d7 */
            {8'h00}, /* 0xd7d6 */
            {8'h00}, /* 0xd7d5 */
            {8'h00}, /* 0xd7d4 */
            {8'h00}, /* 0xd7d3 */
            {8'h00}, /* 0xd7d2 */
            {8'h00}, /* 0xd7d1 */
            {8'h00}, /* 0xd7d0 */
            {8'h00}, /* 0xd7cf */
            {8'h00}, /* 0xd7ce */
            {8'h00}, /* 0xd7cd */
            {8'h00}, /* 0xd7cc */
            {8'h00}, /* 0xd7cb */
            {8'h00}, /* 0xd7ca */
            {8'h00}, /* 0xd7c9 */
            {8'h00}, /* 0xd7c8 */
            {8'h00}, /* 0xd7c7 */
            {8'h00}, /* 0xd7c6 */
            {8'h00}, /* 0xd7c5 */
            {8'h00}, /* 0xd7c4 */
            {8'h00}, /* 0xd7c3 */
            {8'h00}, /* 0xd7c2 */
            {8'h00}, /* 0xd7c1 */
            {8'h00}, /* 0xd7c0 */
            {8'h00}, /* 0xd7bf */
            {8'h00}, /* 0xd7be */
            {8'h00}, /* 0xd7bd */
            {8'h00}, /* 0xd7bc */
            {8'h00}, /* 0xd7bb */
            {8'h00}, /* 0xd7ba */
            {8'h00}, /* 0xd7b9 */
            {8'h00}, /* 0xd7b8 */
            {8'h00}, /* 0xd7b7 */
            {8'h00}, /* 0xd7b6 */
            {8'h00}, /* 0xd7b5 */
            {8'h00}, /* 0xd7b4 */
            {8'h00}, /* 0xd7b3 */
            {8'h00}, /* 0xd7b2 */
            {8'h00}, /* 0xd7b1 */
            {8'h00}, /* 0xd7b0 */
            {8'h00}, /* 0xd7af */
            {8'h00}, /* 0xd7ae */
            {8'h00}, /* 0xd7ad */
            {8'h00}, /* 0xd7ac */
            {8'h00}, /* 0xd7ab */
            {8'h00}, /* 0xd7aa */
            {8'h00}, /* 0xd7a9 */
            {8'h00}, /* 0xd7a8 */
            {8'h00}, /* 0xd7a7 */
            {8'h00}, /* 0xd7a6 */
            {8'h00}, /* 0xd7a5 */
            {8'h00}, /* 0xd7a4 */
            {8'h00}, /* 0xd7a3 */
            {8'h00}, /* 0xd7a2 */
            {8'h00}, /* 0xd7a1 */
            {8'h00}, /* 0xd7a0 */
            {8'h00}, /* 0xd79f */
            {8'h00}, /* 0xd79e */
            {8'h00}, /* 0xd79d */
            {8'h00}, /* 0xd79c */
            {8'h00}, /* 0xd79b */
            {8'h00}, /* 0xd79a */
            {8'h00}, /* 0xd799 */
            {8'h00}, /* 0xd798 */
            {8'h00}, /* 0xd797 */
            {8'h00}, /* 0xd796 */
            {8'h00}, /* 0xd795 */
            {8'h00}, /* 0xd794 */
            {8'h00}, /* 0xd793 */
            {8'h00}, /* 0xd792 */
            {8'h00}, /* 0xd791 */
            {8'h00}, /* 0xd790 */
            {8'h00}, /* 0xd78f */
            {8'h00}, /* 0xd78e */
            {8'h00}, /* 0xd78d */
            {8'h00}, /* 0xd78c */
            {8'h00}, /* 0xd78b */
            {8'h00}, /* 0xd78a */
            {8'h00}, /* 0xd789 */
            {8'h00}, /* 0xd788 */
            {8'h00}, /* 0xd787 */
            {8'h00}, /* 0xd786 */
            {8'h00}, /* 0xd785 */
            {8'h00}, /* 0xd784 */
            {8'h00}, /* 0xd783 */
            {8'h00}, /* 0xd782 */
            {8'h00}, /* 0xd781 */
            {8'h00}, /* 0xd780 */
            {8'h00}, /* 0xd77f */
            {8'h00}, /* 0xd77e */
            {8'h00}, /* 0xd77d */
            {8'h00}, /* 0xd77c */
            {8'h00}, /* 0xd77b */
            {8'h00}, /* 0xd77a */
            {8'h00}, /* 0xd779 */
            {8'h00}, /* 0xd778 */
            {8'h00}, /* 0xd777 */
            {8'h00}, /* 0xd776 */
            {8'h00}, /* 0xd775 */
            {8'h00}, /* 0xd774 */
            {8'h00}, /* 0xd773 */
            {8'h00}, /* 0xd772 */
            {8'h00}, /* 0xd771 */
            {8'h00}, /* 0xd770 */
            {8'h00}, /* 0xd76f */
            {8'h00}, /* 0xd76e */
            {8'h00}, /* 0xd76d */
            {8'h00}, /* 0xd76c */
            {8'h00}, /* 0xd76b */
            {8'h00}, /* 0xd76a */
            {8'h00}, /* 0xd769 */
            {8'h00}, /* 0xd768 */
            {8'h00}, /* 0xd767 */
            {8'h00}, /* 0xd766 */
            {8'h00}, /* 0xd765 */
            {8'h00}, /* 0xd764 */
            {8'h00}, /* 0xd763 */
            {8'h00}, /* 0xd762 */
            {8'h00}, /* 0xd761 */
            {8'h00}, /* 0xd760 */
            {8'h00}, /* 0xd75f */
            {8'h00}, /* 0xd75e */
            {8'h00}, /* 0xd75d */
            {8'h00}, /* 0xd75c */
            {8'h00}, /* 0xd75b */
            {8'h00}, /* 0xd75a */
            {8'h00}, /* 0xd759 */
            {8'h00}, /* 0xd758 */
            {8'h00}, /* 0xd757 */
            {8'h00}, /* 0xd756 */
            {8'h00}, /* 0xd755 */
            {8'h00}, /* 0xd754 */
            {8'h00}, /* 0xd753 */
            {8'h00}, /* 0xd752 */
            {8'h00}, /* 0xd751 */
            {8'h00}, /* 0xd750 */
            {8'h00}, /* 0xd74f */
            {8'h00}, /* 0xd74e */
            {8'h00}, /* 0xd74d */
            {8'h00}, /* 0xd74c */
            {8'h00}, /* 0xd74b */
            {8'h00}, /* 0xd74a */
            {8'h00}, /* 0xd749 */
            {8'h00}, /* 0xd748 */
            {8'h00}, /* 0xd747 */
            {8'h00}, /* 0xd746 */
            {8'h00}, /* 0xd745 */
            {8'h00}, /* 0xd744 */
            {8'h00}, /* 0xd743 */
            {8'h00}, /* 0xd742 */
            {8'h00}, /* 0xd741 */
            {8'h00}, /* 0xd740 */
            {8'h00}, /* 0xd73f */
            {8'h00}, /* 0xd73e */
            {8'h00}, /* 0xd73d */
            {8'h00}, /* 0xd73c */
            {8'h00}, /* 0xd73b */
            {8'h00}, /* 0xd73a */
            {8'h00}, /* 0xd739 */
            {8'h00}, /* 0xd738 */
            {8'h00}, /* 0xd737 */
            {8'h00}, /* 0xd736 */
            {8'h00}, /* 0xd735 */
            {8'h00}, /* 0xd734 */
            {8'h00}, /* 0xd733 */
            {8'h00}, /* 0xd732 */
            {8'h00}, /* 0xd731 */
            {8'h00}, /* 0xd730 */
            {8'h00}, /* 0xd72f */
            {8'h00}, /* 0xd72e */
            {8'h00}, /* 0xd72d */
            {8'h00}, /* 0xd72c */
            {8'h00}, /* 0xd72b */
            {8'h00}, /* 0xd72a */
            {8'h00}, /* 0xd729 */
            {8'h00}, /* 0xd728 */
            {8'h00}, /* 0xd727 */
            {8'h00}, /* 0xd726 */
            {8'h00}, /* 0xd725 */
            {8'h00}, /* 0xd724 */
            {8'h00}, /* 0xd723 */
            {8'h00}, /* 0xd722 */
            {8'h00}, /* 0xd721 */
            {8'h00}, /* 0xd720 */
            {8'h00}, /* 0xd71f */
            {8'h00}, /* 0xd71e */
            {8'h00}, /* 0xd71d */
            {8'h00}, /* 0xd71c */
            {8'h00}, /* 0xd71b */
            {8'h00}, /* 0xd71a */
            {8'h00}, /* 0xd719 */
            {8'h00}, /* 0xd718 */
            {8'h00}, /* 0xd717 */
            {8'h00}, /* 0xd716 */
            {8'h00}, /* 0xd715 */
            {8'h00}, /* 0xd714 */
            {8'h00}, /* 0xd713 */
            {8'h00}, /* 0xd712 */
            {8'h00}, /* 0xd711 */
            {8'h00}, /* 0xd710 */
            {8'h00}, /* 0xd70f */
            {8'h00}, /* 0xd70e */
            {8'h00}, /* 0xd70d */
            {8'h00}, /* 0xd70c */
            {8'h00}, /* 0xd70b */
            {8'h00}, /* 0xd70a */
            {8'h00}, /* 0xd709 */
            {8'h00}, /* 0xd708 */
            {8'h00}, /* 0xd707 */
            {8'h00}, /* 0xd706 */
            {8'h00}, /* 0xd705 */
            {8'h00}, /* 0xd704 */
            {8'h00}, /* 0xd703 */
            {8'h00}, /* 0xd702 */
            {8'h00}, /* 0xd701 */
            {8'h00}, /* 0xd700 */
            {8'h00}, /* 0xd6ff */
            {8'h00}, /* 0xd6fe */
            {8'h00}, /* 0xd6fd */
            {8'h00}, /* 0xd6fc */
            {8'h00}, /* 0xd6fb */
            {8'h00}, /* 0xd6fa */
            {8'h00}, /* 0xd6f9 */
            {8'h00}, /* 0xd6f8 */
            {8'h00}, /* 0xd6f7 */
            {8'h00}, /* 0xd6f6 */
            {8'h00}, /* 0xd6f5 */
            {8'h00}, /* 0xd6f4 */
            {8'h00}, /* 0xd6f3 */
            {8'h00}, /* 0xd6f2 */
            {8'h00}, /* 0xd6f1 */
            {8'h00}, /* 0xd6f0 */
            {8'h00}, /* 0xd6ef */
            {8'h00}, /* 0xd6ee */
            {8'h00}, /* 0xd6ed */
            {8'h00}, /* 0xd6ec */
            {8'h00}, /* 0xd6eb */
            {8'h00}, /* 0xd6ea */
            {8'h00}, /* 0xd6e9 */
            {8'h00}, /* 0xd6e8 */
            {8'h00}, /* 0xd6e7 */
            {8'h00}, /* 0xd6e6 */
            {8'h00}, /* 0xd6e5 */
            {8'h00}, /* 0xd6e4 */
            {8'h00}, /* 0xd6e3 */
            {8'h00}, /* 0xd6e2 */
            {8'h00}, /* 0xd6e1 */
            {8'h00}, /* 0xd6e0 */
            {8'h00}, /* 0xd6df */
            {8'h00}, /* 0xd6de */
            {8'h00}, /* 0xd6dd */
            {8'h00}, /* 0xd6dc */
            {8'h00}, /* 0xd6db */
            {8'h00}, /* 0xd6da */
            {8'h00}, /* 0xd6d9 */
            {8'h00}, /* 0xd6d8 */
            {8'h00}, /* 0xd6d7 */
            {8'h00}, /* 0xd6d6 */
            {8'h00}, /* 0xd6d5 */
            {8'h00}, /* 0xd6d4 */
            {8'h00}, /* 0xd6d3 */
            {8'h00}, /* 0xd6d2 */
            {8'h00}, /* 0xd6d1 */
            {8'h00}, /* 0xd6d0 */
            {8'h00}, /* 0xd6cf */
            {8'h00}, /* 0xd6ce */
            {8'h00}, /* 0xd6cd */
            {8'h00}, /* 0xd6cc */
            {8'h00}, /* 0xd6cb */
            {8'h00}, /* 0xd6ca */
            {8'h00}, /* 0xd6c9 */
            {8'h00}, /* 0xd6c8 */
            {8'h00}, /* 0xd6c7 */
            {8'h00}, /* 0xd6c6 */
            {8'h00}, /* 0xd6c5 */
            {8'h00}, /* 0xd6c4 */
            {8'h00}, /* 0xd6c3 */
            {8'h00}, /* 0xd6c2 */
            {8'h00}, /* 0xd6c1 */
            {8'h00}, /* 0xd6c0 */
            {8'h00}, /* 0xd6bf */
            {8'h00}, /* 0xd6be */
            {8'h00}, /* 0xd6bd */
            {8'h00}, /* 0xd6bc */
            {8'h00}, /* 0xd6bb */
            {8'h00}, /* 0xd6ba */
            {8'h00}, /* 0xd6b9 */
            {8'h00}, /* 0xd6b8 */
            {8'h00}, /* 0xd6b7 */
            {8'h00}, /* 0xd6b6 */
            {8'h00}, /* 0xd6b5 */
            {8'h00}, /* 0xd6b4 */
            {8'h00}, /* 0xd6b3 */
            {8'h00}, /* 0xd6b2 */
            {8'h00}, /* 0xd6b1 */
            {8'h00}, /* 0xd6b0 */
            {8'h00}, /* 0xd6af */
            {8'h00}, /* 0xd6ae */
            {8'h00}, /* 0xd6ad */
            {8'h00}, /* 0xd6ac */
            {8'h00}, /* 0xd6ab */
            {8'h00}, /* 0xd6aa */
            {8'h00}, /* 0xd6a9 */
            {8'h00}, /* 0xd6a8 */
            {8'h00}, /* 0xd6a7 */
            {8'h00}, /* 0xd6a6 */
            {8'h00}, /* 0xd6a5 */
            {8'h00}, /* 0xd6a4 */
            {8'h00}, /* 0xd6a3 */
            {8'h00}, /* 0xd6a2 */
            {8'h00}, /* 0xd6a1 */
            {8'h00}, /* 0xd6a0 */
            {8'h00}, /* 0xd69f */
            {8'h00}, /* 0xd69e */
            {8'h00}, /* 0xd69d */
            {8'h00}, /* 0xd69c */
            {8'h00}, /* 0xd69b */
            {8'h00}, /* 0xd69a */
            {8'h00}, /* 0xd699 */
            {8'h00}, /* 0xd698 */
            {8'h00}, /* 0xd697 */
            {8'h00}, /* 0xd696 */
            {8'h00}, /* 0xd695 */
            {8'h00}, /* 0xd694 */
            {8'h00}, /* 0xd693 */
            {8'h00}, /* 0xd692 */
            {8'h00}, /* 0xd691 */
            {8'h00}, /* 0xd690 */
            {8'h00}, /* 0xd68f */
            {8'h00}, /* 0xd68e */
            {8'h00}, /* 0xd68d */
            {8'h00}, /* 0xd68c */
            {8'h00}, /* 0xd68b */
            {8'h00}, /* 0xd68a */
            {8'h00}, /* 0xd689 */
            {8'h00}, /* 0xd688 */
            {8'h00}, /* 0xd687 */
            {8'h00}, /* 0xd686 */
            {8'h00}, /* 0xd685 */
            {8'h00}, /* 0xd684 */
            {8'h00}, /* 0xd683 */
            {8'h00}, /* 0xd682 */
            {8'h00}, /* 0xd681 */
            {8'h00}, /* 0xd680 */
            {8'h00}, /* 0xd67f */
            {8'h00}, /* 0xd67e */
            {8'h00}, /* 0xd67d */
            {8'h00}, /* 0xd67c */
            {8'h00}, /* 0xd67b */
            {8'h00}, /* 0xd67a */
            {8'h00}, /* 0xd679 */
            {8'h00}, /* 0xd678 */
            {8'h00}, /* 0xd677 */
            {8'h00}, /* 0xd676 */
            {8'h00}, /* 0xd675 */
            {8'h00}, /* 0xd674 */
            {8'h00}, /* 0xd673 */
            {8'h00}, /* 0xd672 */
            {8'h00}, /* 0xd671 */
            {8'h00}, /* 0xd670 */
            {8'h00}, /* 0xd66f */
            {8'h00}, /* 0xd66e */
            {8'h00}, /* 0xd66d */
            {8'h00}, /* 0xd66c */
            {8'h00}, /* 0xd66b */
            {8'h00}, /* 0xd66a */
            {8'h00}, /* 0xd669 */
            {8'h00}, /* 0xd668 */
            {8'h00}, /* 0xd667 */
            {8'h00}, /* 0xd666 */
            {8'h00}, /* 0xd665 */
            {8'h00}, /* 0xd664 */
            {8'h00}, /* 0xd663 */
            {8'h00}, /* 0xd662 */
            {8'h00}, /* 0xd661 */
            {8'h00}, /* 0xd660 */
            {8'h00}, /* 0xd65f */
            {8'h00}, /* 0xd65e */
            {8'h00}, /* 0xd65d */
            {8'h00}, /* 0xd65c */
            {8'h00}, /* 0xd65b */
            {8'h00}, /* 0xd65a */
            {8'h00}, /* 0xd659 */
            {8'h00}, /* 0xd658 */
            {8'h00}, /* 0xd657 */
            {8'h00}, /* 0xd656 */
            {8'h00}, /* 0xd655 */
            {8'h00}, /* 0xd654 */
            {8'h00}, /* 0xd653 */
            {8'h00}, /* 0xd652 */
            {8'h00}, /* 0xd651 */
            {8'h00}, /* 0xd650 */
            {8'h00}, /* 0xd64f */
            {8'h00}, /* 0xd64e */
            {8'h00}, /* 0xd64d */
            {8'h00}, /* 0xd64c */
            {8'h00}, /* 0xd64b */
            {8'h00}, /* 0xd64a */
            {8'h00}, /* 0xd649 */
            {8'h00}, /* 0xd648 */
            {8'h00}, /* 0xd647 */
            {8'h00}, /* 0xd646 */
            {8'h00}, /* 0xd645 */
            {8'h00}, /* 0xd644 */
            {8'h00}, /* 0xd643 */
            {8'h00}, /* 0xd642 */
            {8'h00}, /* 0xd641 */
            {8'h00}, /* 0xd640 */
            {8'h00}, /* 0xd63f */
            {8'h00}, /* 0xd63e */
            {8'h00}, /* 0xd63d */
            {8'h00}, /* 0xd63c */
            {8'h00}, /* 0xd63b */
            {8'h00}, /* 0xd63a */
            {8'h00}, /* 0xd639 */
            {8'h00}, /* 0xd638 */
            {8'h00}, /* 0xd637 */
            {8'h00}, /* 0xd636 */
            {8'h00}, /* 0xd635 */
            {8'h00}, /* 0xd634 */
            {8'h00}, /* 0xd633 */
            {8'h00}, /* 0xd632 */
            {8'h00}, /* 0xd631 */
            {8'h00}, /* 0xd630 */
            {8'h00}, /* 0xd62f */
            {8'h00}, /* 0xd62e */
            {8'h00}, /* 0xd62d */
            {8'h00}, /* 0xd62c */
            {8'h00}, /* 0xd62b */
            {8'h00}, /* 0xd62a */
            {8'h00}, /* 0xd629 */
            {8'h00}, /* 0xd628 */
            {8'h00}, /* 0xd627 */
            {8'h00}, /* 0xd626 */
            {8'h00}, /* 0xd625 */
            {8'h00}, /* 0xd624 */
            {8'h00}, /* 0xd623 */
            {8'h00}, /* 0xd622 */
            {8'h00}, /* 0xd621 */
            {8'h00}, /* 0xd620 */
            {8'h00}, /* 0xd61f */
            {8'h00}, /* 0xd61e */
            {8'h00}, /* 0xd61d */
            {8'h00}, /* 0xd61c */
            {8'h00}, /* 0xd61b */
            {8'h00}, /* 0xd61a */
            {8'h00}, /* 0xd619 */
            {8'h00}, /* 0xd618 */
            {8'h00}, /* 0xd617 */
            {8'h00}, /* 0xd616 */
            {8'h00}, /* 0xd615 */
            {8'h00}, /* 0xd614 */
            {8'h00}, /* 0xd613 */
            {8'h00}, /* 0xd612 */
            {8'h00}, /* 0xd611 */
            {8'h00}, /* 0xd610 */
            {8'h00}, /* 0xd60f */
            {8'h00}, /* 0xd60e */
            {8'h00}, /* 0xd60d */
            {8'h00}, /* 0xd60c */
            {8'h00}, /* 0xd60b */
            {8'h00}, /* 0xd60a */
            {8'h00}, /* 0xd609 */
            {8'h00}, /* 0xd608 */
            {8'h00}, /* 0xd607 */
            {8'h00}, /* 0xd606 */
            {8'h00}, /* 0xd605 */
            {8'h00}, /* 0xd604 */
            {8'h00}, /* 0xd603 */
            {8'h00}, /* 0xd602 */
            {8'h00}, /* 0xd601 */
            {8'h00}, /* 0xd600 */
            {8'h00}, /* 0xd5ff */
            {8'h00}, /* 0xd5fe */
            {8'h00}, /* 0xd5fd */
            {8'h00}, /* 0xd5fc */
            {8'h00}, /* 0xd5fb */
            {8'h00}, /* 0xd5fa */
            {8'h00}, /* 0xd5f9 */
            {8'h00}, /* 0xd5f8 */
            {8'h00}, /* 0xd5f7 */
            {8'h00}, /* 0xd5f6 */
            {8'h00}, /* 0xd5f5 */
            {8'h00}, /* 0xd5f4 */
            {8'h00}, /* 0xd5f3 */
            {8'h00}, /* 0xd5f2 */
            {8'h00}, /* 0xd5f1 */
            {8'h00}, /* 0xd5f0 */
            {8'h00}, /* 0xd5ef */
            {8'h00}, /* 0xd5ee */
            {8'h00}, /* 0xd5ed */
            {8'h00}, /* 0xd5ec */
            {8'h00}, /* 0xd5eb */
            {8'h00}, /* 0xd5ea */
            {8'h00}, /* 0xd5e9 */
            {8'h00}, /* 0xd5e8 */
            {8'h00}, /* 0xd5e7 */
            {8'h00}, /* 0xd5e6 */
            {8'h00}, /* 0xd5e5 */
            {8'h00}, /* 0xd5e4 */
            {8'h00}, /* 0xd5e3 */
            {8'h00}, /* 0xd5e2 */
            {8'h00}, /* 0xd5e1 */
            {8'h00}, /* 0xd5e0 */
            {8'h00}, /* 0xd5df */
            {8'h00}, /* 0xd5de */
            {8'h00}, /* 0xd5dd */
            {8'h00}, /* 0xd5dc */
            {8'h00}, /* 0xd5db */
            {8'h00}, /* 0xd5da */
            {8'h00}, /* 0xd5d9 */
            {8'h00}, /* 0xd5d8 */
            {8'h00}, /* 0xd5d7 */
            {8'h00}, /* 0xd5d6 */
            {8'h00}, /* 0xd5d5 */
            {8'h00}, /* 0xd5d4 */
            {8'h00}, /* 0xd5d3 */
            {8'h00}, /* 0xd5d2 */
            {8'h00}, /* 0xd5d1 */
            {8'h00}, /* 0xd5d0 */
            {8'h00}, /* 0xd5cf */
            {8'h00}, /* 0xd5ce */
            {8'h00}, /* 0xd5cd */
            {8'h00}, /* 0xd5cc */
            {8'h00}, /* 0xd5cb */
            {8'h00}, /* 0xd5ca */
            {8'h00}, /* 0xd5c9 */
            {8'h00}, /* 0xd5c8 */
            {8'h00}, /* 0xd5c7 */
            {8'h00}, /* 0xd5c6 */
            {8'h00}, /* 0xd5c5 */
            {8'h00}, /* 0xd5c4 */
            {8'h00}, /* 0xd5c3 */
            {8'h00}, /* 0xd5c2 */
            {8'h00}, /* 0xd5c1 */
            {8'h00}, /* 0xd5c0 */
            {8'h00}, /* 0xd5bf */
            {8'h00}, /* 0xd5be */
            {8'h00}, /* 0xd5bd */
            {8'h00}, /* 0xd5bc */
            {8'h00}, /* 0xd5bb */
            {8'h00}, /* 0xd5ba */
            {8'h00}, /* 0xd5b9 */
            {8'h00}, /* 0xd5b8 */
            {8'h00}, /* 0xd5b7 */
            {8'h00}, /* 0xd5b6 */
            {8'h00}, /* 0xd5b5 */
            {8'h00}, /* 0xd5b4 */
            {8'h00}, /* 0xd5b3 */
            {8'h00}, /* 0xd5b2 */
            {8'h00}, /* 0xd5b1 */
            {8'h00}, /* 0xd5b0 */
            {8'h00}, /* 0xd5af */
            {8'h00}, /* 0xd5ae */
            {8'h00}, /* 0xd5ad */
            {8'h00}, /* 0xd5ac */
            {8'h00}, /* 0xd5ab */
            {8'h00}, /* 0xd5aa */
            {8'h00}, /* 0xd5a9 */
            {8'h00}, /* 0xd5a8 */
            {8'h00}, /* 0xd5a7 */
            {8'h00}, /* 0xd5a6 */
            {8'h00}, /* 0xd5a5 */
            {8'h00}, /* 0xd5a4 */
            {8'h00}, /* 0xd5a3 */
            {8'h00}, /* 0xd5a2 */
            {8'h00}, /* 0xd5a1 */
            {8'h00}, /* 0xd5a0 */
            {8'h00}, /* 0xd59f */
            {8'h00}, /* 0xd59e */
            {8'h00}, /* 0xd59d */
            {8'h00}, /* 0xd59c */
            {8'h00}, /* 0xd59b */
            {8'h00}, /* 0xd59a */
            {8'h00}, /* 0xd599 */
            {8'h00}, /* 0xd598 */
            {8'h00}, /* 0xd597 */
            {8'h00}, /* 0xd596 */
            {8'h00}, /* 0xd595 */
            {8'h00}, /* 0xd594 */
            {8'h00}, /* 0xd593 */
            {8'h00}, /* 0xd592 */
            {8'h00}, /* 0xd591 */
            {8'h00}, /* 0xd590 */
            {8'h00}, /* 0xd58f */
            {8'h00}, /* 0xd58e */
            {8'h00}, /* 0xd58d */
            {8'h00}, /* 0xd58c */
            {8'h00}, /* 0xd58b */
            {8'h00}, /* 0xd58a */
            {8'h00}, /* 0xd589 */
            {8'h00}, /* 0xd588 */
            {8'h00}, /* 0xd587 */
            {8'h00}, /* 0xd586 */
            {8'h00}, /* 0xd585 */
            {8'h00}, /* 0xd584 */
            {8'h00}, /* 0xd583 */
            {8'h00}, /* 0xd582 */
            {8'h00}, /* 0xd581 */
            {8'h00}, /* 0xd580 */
            {8'h00}, /* 0xd57f */
            {8'h00}, /* 0xd57e */
            {8'h00}, /* 0xd57d */
            {8'h00}, /* 0xd57c */
            {8'h00}, /* 0xd57b */
            {8'h00}, /* 0xd57a */
            {8'h00}, /* 0xd579 */
            {8'h00}, /* 0xd578 */
            {8'h00}, /* 0xd577 */
            {8'h00}, /* 0xd576 */
            {8'h00}, /* 0xd575 */
            {8'h00}, /* 0xd574 */
            {8'h00}, /* 0xd573 */
            {8'h00}, /* 0xd572 */
            {8'h00}, /* 0xd571 */
            {8'h00}, /* 0xd570 */
            {8'h00}, /* 0xd56f */
            {8'h00}, /* 0xd56e */
            {8'h00}, /* 0xd56d */
            {8'h00}, /* 0xd56c */
            {8'h00}, /* 0xd56b */
            {8'h00}, /* 0xd56a */
            {8'h00}, /* 0xd569 */
            {8'h00}, /* 0xd568 */
            {8'h00}, /* 0xd567 */
            {8'h00}, /* 0xd566 */
            {8'h00}, /* 0xd565 */
            {8'h00}, /* 0xd564 */
            {8'h00}, /* 0xd563 */
            {8'h00}, /* 0xd562 */
            {8'h00}, /* 0xd561 */
            {8'h00}, /* 0xd560 */
            {8'h00}, /* 0xd55f */
            {8'h00}, /* 0xd55e */
            {8'h00}, /* 0xd55d */
            {8'h00}, /* 0xd55c */
            {8'h00}, /* 0xd55b */
            {8'h00}, /* 0xd55a */
            {8'h00}, /* 0xd559 */
            {8'h00}, /* 0xd558 */
            {8'h00}, /* 0xd557 */
            {8'h00}, /* 0xd556 */
            {8'h00}, /* 0xd555 */
            {8'h00}, /* 0xd554 */
            {8'h00}, /* 0xd553 */
            {8'h00}, /* 0xd552 */
            {8'h00}, /* 0xd551 */
            {8'h00}, /* 0xd550 */
            {8'h00}, /* 0xd54f */
            {8'h00}, /* 0xd54e */
            {8'h00}, /* 0xd54d */
            {8'h00}, /* 0xd54c */
            {8'h00}, /* 0xd54b */
            {8'h00}, /* 0xd54a */
            {8'h00}, /* 0xd549 */
            {8'h00}, /* 0xd548 */
            {8'h00}, /* 0xd547 */
            {8'h00}, /* 0xd546 */
            {8'h00}, /* 0xd545 */
            {8'h00}, /* 0xd544 */
            {8'h00}, /* 0xd543 */
            {8'h00}, /* 0xd542 */
            {8'h00}, /* 0xd541 */
            {8'h00}, /* 0xd540 */
            {8'h00}, /* 0xd53f */
            {8'h00}, /* 0xd53e */
            {8'h00}, /* 0xd53d */
            {8'h00}, /* 0xd53c */
            {8'h00}, /* 0xd53b */
            {8'h00}, /* 0xd53a */
            {8'h00}, /* 0xd539 */
            {8'h00}, /* 0xd538 */
            {8'h00}, /* 0xd537 */
            {8'h00}, /* 0xd536 */
            {8'h00}, /* 0xd535 */
            {8'h00}, /* 0xd534 */
            {8'h00}, /* 0xd533 */
            {8'h00}, /* 0xd532 */
            {8'h00}, /* 0xd531 */
            {8'h00}, /* 0xd530 */
            {8'h00}, /* 0xd52f */
            {8'h00}, /* 0xd52e */
            {8'h00}, /* 0xd52d */
            {8'h00}, /* 0xd52c */
            {8'h00}, /* 0xd52b */
            {8'h00}, /* 0xd52a */
            {8'h00}, /* 0xd529 */
            {8'h00}, /* 0xd528 */
            {8'h00}, /* 0xd527 */
            {8'h00}, /* 0xd526 */
            {8'h00}, /* 0xd525 */
            {8'h00}, /* 0xd524 */
            {8'h00}, /* 0xd523 */
            {8'h00}, /* 0xd522 */
            {8'h00}, /* 0xd521 */
            {8'h00}, /* 0xd520 */
            {8'h00}, /* 0xd51f */
            {8'h00}, /* 0xd51e */
            {8'h00}, /* 0xd51d */
            {8'h00}, /* 0xd51c */
            {8'h00}, /* 0xd51b */
            {8'h00}, /* 0xd51a */
            {8'h00}, /* 0xd519 */
            {8'h00}, /* 0xd518 */
            {8'h00}, /* 0xd517 */
            {8'h00}, /* 0xd516 */
            {8'h00}, /* 0xd515 */
            {8'h00}, /* 0xd514 */
            {8'h00}, /* 0xd513 */
            {8'h00}, /* 0xd512 */
            {8'h00}, /* 0xd511 */
            {8'h00}, /* 0xd510 */
            {8'h00}, /* 0xd50f */
            {8'h00}, /* 0xd50e */
            {8'h00}, /* 0xd50d */
            {8'h00}, /* 0xd50c */
            {8'h00}, /* 0xd50b */
            {8'h00}, /* 0xd50a */
            {8'h00}, /* 0xd509 */
            {8'h00}, /* 0xd508 */
            {8'h00}, /* 0xd507 */
            {8'h00}, /* 0xd506 */
            {8'h00}, /* 0xd505 */
            {8'h00}, /* 0xd504 */
            {8'h00}, /* 0xd503 */
            {8'h00}, /* 0xd502 */
            {8'h00}, /* 0xd501 */
            {8'h00}, /* 0xd500 */
            {8'h00}, /* 0xd4ff */
            {8'h00}, /* 0xd4fe */
            {8'h00}, /* 0xd4fd */
            {8'h00}, /* 0xd4fc */
            {8'h00}, /* 0xd4fb */
            {8'h00}, /* 0xd4fa */
            {8'h00}, /* 0xd4f9 */
            {8'h00}, /* 0xd4f8 */
            {8'h00}, /* 0xd4f7 */
            {8'h00}, /* 0xd4f6 */
            {8'h00}, /* 0xd4f5 */
            {8'h00}, /* 0xd4f4 */
            {8'h00}, /* 0xd4f3 */
            {8'h00}, /* 0xd4f2 */
            {8'h00}, /* 0xd4f1 */
            {8'h00}, /* 0xd4f0 */
            {8'h00}, /* 0xd4ef */
            {8'h00}, /* 0xd4ee */
            {8'h00}, /* 0xd4ed */
            {8'h00}, /* 0xd4ec */
            {8'h00}, /* 0xd4eb */
            {8'h00}, /* 0xd4ea */
            {8'h00}, /* 0xd4e9 */
            {8'h00}, /* 0xd4e8 */
            {8'h00}, /* 0xd4e7 */
            {8'h00}, /* 0xd4e6 */
            {8'h00}, /* 0xd4e5 */
            {8'h00}, /* 0xd4e4 */
            {8'h00}, /* 0xd4e3 */
            {8'h00}, /* 0xd4e2 */
            {8'h00}, /* 0xd4e1 */
            {8'h00}, /* 0xd4e0 */
            {8'h00}, /* 0xd4df */
            {8'h00}, /* 0xd4de */
            {8'h00}, /* 0xd4dd */
            {8'h00}, /* 0xd4dc */
            {8'h00}, /* 0xd4db */
            {8'h00}, /* 0xd4da */
            {8'h00}, /* 0xd4d9 */
            {8'h00}, /* 0xd4d8 */
            {8'h00}, /* 0xd4d7 */
            {8'h00}, /* 0xd4d6 */
            {8'h00}, /* 0xd4d5 */
            {8'h00}, /* 0xd4d4 */
            {8'h00}, /* 0xd4d3 */
            {8'h00}, /* 0xd4d2 */
            {8'h00}, /* 0xd4d1 */
            {8'h00}, /* 0xd4d0 */
            {8'h00}, /* 0xd4cf */
            {8'h00}, /* 0xd4ce */
            {8'h00}, /* 0xd4cd */
            {8'h00}, /* 0xd4cc */
            {8'h00}, /* 0xd4cb */
            {8'h00}, /* 0xd4ca */
            {8'h00}, /* 0xd4c9 */
            {8'h00}, /* 0xd4c8 */
            {8'h00}, /* 0xd4c7 */
            {8'h00}, /* 0xd4c6 */
            {8'h00}, /* 0xd4c5 */
            {8'h00}, /* 0xd4c4 */
            {8'h00}, /* 0xd4c3 */
            {8'h00}, /* 0xd4c2 */
            {8'h00}, /* 0xd4c1 */
            {8'h00}, /* 0xd4c0 */
            {8'h00}, /* 0xd4bf */
            {8'h00}, /* 0xd4be */
            {8'h00}, /* 0xd4bd */
            {8'h00}, /* 0xd4bc */
            {8'h00}, /* 0xd4bb */
            {8'h00}, /* 0xd4ba */
            {8'h00}, /* 0xd4b9 */
            {8'h00}, /* 0xd4b8 */
            {8'h00}, /* 0xd4b7 */
            {8'h00}, /* 0xd4b6 */
            {8'h00}, /* 0xd4b5 */
            {8'h00}, /* 0xd4b4 */
            {8'h00}, /* 0xd4b3 */
            {8'h00}, /* 0xd4b2 */
            {8'h00}, /* 0xd4b1 */
            {8'h00}, /* 0xd4b0 */
            {8'h00}, /* 0xd4af */
            {8'h00}, /* 0xd4ae */
            {8'h00}, /* 0xd4ad */
            {8'h00}, /* 0xd4ac */
            {8'h00}, /* 0xd4ab */
            {8'h00}, /* 0xd4aa */
            {8'h00}, /* 0xd4a9 */
            {8'h00}, /* 0xd4a8 */
            {8'h00}, /* 0xd4a7 */
            {8'h00}, /* 0xd4a6 */
            {8'h00}, /* 0xd4a5 */
            {8'h00}, /* 0xd4a4 */
            {8'h00}, /* 0xd4a3 */
            {8'h00}, /* 0xd4a2 */
            {8'h00}, /* 0xd4a1 */
            {8'h00}, /* 0xd4a0 */
            {8'h00}, /* 0xd49f */
            {8'h00}, /* 0xd49e */
            {8'h00}, /* 0xd49d */
            {8'h00}, /* 0xd49c */
            {8'h00}, /* 0xd49b */
            {8'h00}, /* 0xd49a */
            {8'h00}, /* 0xd499 */
            {8'h00}, /* 0xd498 */
            {8'h00}, /* 0xd497 */
            {8'h00}, /* 0xd496 */
            {8'h00}, /* 0xd495 */
            {8'h00}, /* 0xd494 */
            {8'h00}, /* 0xd493 */
            {8'h00}, /* 0xd492 */
            {8'h00}, /* 0xd491 */
            {8'h00}, /* 0xd490 */
            {8'h00}, /* 0xd48f */
            {8'h00}, /* 0xd48e */
            {8'h00}, /* 0xd48d */
            {8'h00}, /* 0xd48c */
            {8'h00}, /* 0xd48b */
            {8'h00}, /* 0xd48a */
            {8'h00}, /* 0xd489 */
            {8'h00}, /* 0xd488 */
            {8'h00}, /* 0xd487 */
            {8'h00}, /* 0xd486 */
            {8'h00}, /* 0xd485 */
            {8'h00}, /* 0xd484 */
            {8'h00}, /* 0xd483 */
            {8'h00}, /* 0xd482 */
            {8'h00}, /* 0xd481 */
            {8'h00}, /* 0xd480 */
            {8'h00}, /* 0xd47f */
            {8'h00}, /* 0xd47e */
            {8'h00}, /* 0xd47d */
            {8'h00}, /* 0xd47c */
            {8'h00}, /* 0xd47b */
            {8'h00}, /* 0xd47a */
            {8'h00}, /* 0xd479 */
            {8'h00}, /* 0xd478 */
            {8'h00}, /* 0xd477 */
            {8'h00}, /* 0xd476 */
            {8'h00}, /* 0xd475 */
            {8'h00}, /* 0xd474 */
            {8'h00}, /* 0xd473 */
            {8'h00}, /* 0xd472 */
            {8'h00}, /* 0xd471 */
            {8'h00}, /* 0xd470 */
            {8'h00}, /* 0xd46f */
            {8'h00}, /* 0xd46e */
            {8'h00}, /* 0xd46d */
            {8'h00}, /* 0xd46c */
            {8'h00}, /* 0xd46b */
            {8'h00}, /* 0xd46a */
            {8'h00}, /* 0xd469 */
            {8'h00}, /* 0xd468 */
            {8'h00}, /* 0xd467 */
            {8'h00}, /* 0xd466 */
            {8'h00}, /* 0xd465 */
            {8'h00}, /* 0xd464 */
            {8'h00}, /* 0xd463 */
            {8'h00}, /* 0xd462 */
            {8'h00}, /* 0xd461 */
            {8'h00}, /* 0xd460 */
            {8'h00}, /* 0xd45f */
            {8'h00}, /* 0xd45e */
            {8'h00}, /* 0xd45d */
            {8'h00}, /* 0xd45c */
            {8'h00}, /* 0xd45b */
            {8'h00}, /* 0xd45a */
            {8'h00}, /* 0xd459 */
            {8'h00}, /* 0xd458 */
            {8'h00}, /* 0xd457 */
            {8'h00}, /* 0xd456 */
            {8'h00}, /* 0xd455 */
            {8'h00}, /* 0xd454 */
            {8'h00}, /* 0xd453 */
            {8'h00}, /* 0xd452 */
            {8'h00}, /* 0xd451 */
            {8'h00}, /* 0xd450 */
            {8'h00}, /* 0xd44f */
            {8'h00}, /* 0xd44e */
            {8'h00}, /* 0xd44d */
            {8'h00}, /* 0xd44c */
            {8'h00}, /* 0xd44b */
            {8'h00}, /* 0xd44a */
            {8'h00}, /* 0xd449 */
            {8'h00}, /* 0xd448 */
            {8'h00}, /* 0xd447 */
            {8'h00}, /* 0xd446 */
            {8'h00}, /* 0xd445 */
            {8'h00}, /* 0xd444 */
            {8'h00}, /* 0xd443 */
            {8'h00}, /* 0xd442 */
            {8'h00}, /* 0xd441 */
            {8'h00}, /* 0xd440 */
            {8'h00}, /* 0xd43f */
            {8'h00}, /* 0xd43e */
            {8'h00}, /* 0xd43d */
            {8'h00}, /* 0xd43c */
            {8'h00}, /* 0xd43b */
            {8'h00}, /* 0xd43a */
            {8'h00}, /* 0xd439 */
            {8'h00}, /* 0xd438 */
            {8'h00}, /* 0xd437 */
            {8'h00}, /* 0xd436 */
            {8'h00}, /* 0xd435 */
            {8'h00}, /* 0xd434 */
            {8'h00}, /* 0xd433 */
            {8'h00}, /* 0xd432 */
            {8'h00}, /* 0xd431 */
            {8'h00}, /* 0xd430 */
            {8'h00}, /* 0xd42f */
            {8'h00}, /* 0xd42e */
            {8'h00}, /* 0xd42d */
            {8'h00}, /* 0xd42c */
            {8'h00}, /* 0xd42b */
            {8'h00}, /* 0xd42a */
            {8'h00}, /* 0xd429 */
            {8'h00}, /* 0xd428 */
            {8'h00}, /* 0xd427 */
            {8'h00}, /* 0xd426 */
            {8'h00}, /* 0xd425 */
            {8'h00}, /* 0xd424 */
            {8'h00}, /* 0xd423 */
            {8'h00}, /* 0xd422 */
            {8'h00}, /* 0xd421 */
            {8'h00}, /* 0xd420 */
            {8'h00}, /* 0xd41f */
            {8'h00}, /* 0xd41e */
            {8'h00}, /* 0xd41d */
            {8'h00}, /* 0xd41c */
            {8'h00}, /* 0xd41b */
            {8'h00}, /* 0xd41a */
            {8'h00}, /* 0xd419 */
            {8'h00}, /* 0xd418 */
            {8'h00}, /* 0xd417 */
            {8'h00}, /* 0xd416 */
            {8'h00}, /* 0xd415 */
            {8'h00}, /* 0xd414 */
            {8'h00}, /* 0xd413 */
            {8'h00}, /* 0xd412 */
            {8'h00}, /* 0xd411 */
            {8'h00}, /* 0xd410 */
            {8'h00}, /* 0xd40f */
            {8'h00}, /* 0xd40e */
            {8'h00}, /* 0xd40d */
            {8'h00}, /* 0xd40c */
            {8'h00}, /* 0xd40b */
            {8'h00}, /* 0xd40a */
            {8'h00}, /* 0xd409 */
            {8'h00}, /* 0xd408 */
            {8'h00}, /* 0xd407 */
            {8'h00}, /* 0xd406 */
            {8'h00}, /* 0xd405 */
            {8'h00}, /* 0xd404 */
            {8'h00}, /* 0xd403 */
            {8'h00}, /* 0xd402 */
            {8'h00}, /* 0xd401 */
            {8'h00}, /* 0xd400 */
            {8'h00}, /* 0xd3ff */
            {8'h00}, /* 0xd3fe */
            {8'h00}, /* 0xd3fd */
            {8'h00}, /* 0xd3fc */
            {8'h00}, /* 0xd3fb */
            {8'h00}, /* 0xd3fa */
            {8'h00}, /* 0xd3f9 */
            {8'h00}, /* 0xd3f8 */
            {8'h00}, /* 0xd3f7 */
            {8'h00}, /* 0xd3f6 */
            {8'h00}, /* 0xd3f5 */
            {8'h00}, /* 0xd3f4 */
            {8'h00}, /* 0xd3f3 */
            {8'h00}, /* 0xd3f2 */
            {8'h00}, /* 0xd3f1 */
            {8'h00}, /* 0xd3f0 */
            {8'h00}, /* 0xd3ef */
            {8'h00}, /* 0xd3ee */
            {8'h00}, /* 0xd3ed */
            {8'h00}, /* 0xd3ec */
            {8'h00}, /* 0xd3eb */
            {8'h00}, /* 0xd3ea */
            {8'h00}, /* 0xd3e9 */
            {8'h00}, /* 0xd3e8 */
            {8'h00}, /* 0xd3e7 */
            {8'h00}, /* 0xd3e6 */
            {8'h00}, /* 0xd3e5 */
            {8'h00}, /* 0xd3e4 */
            {8'h00}, /* 0xd3e3 */
            {8'h00}, /* 0xd3e2 */
            {8'h00}, /* 0xd3e1 */
            {8'h00}, /* 0xd3e0 */
            {8'h00}, /* 0xd3df */
            {8'h00}, /* 0xd3de */
            {8'h00}, /* 0xd3dd */
            {8'h00}, /* 0xd3dc */
            {8'h00}, /* 0xd3db */
            {8'h00}, /* 0xd3da */
            {8'h00}, /* 0xd3d9 */
            {8'h00}, /* 0xd3d8 */
            {8'h00}, /* 0xd3d7 */
            {8'h00}, /* 0xd3d6 */
            {8'h00}, /* 0xd3d5 */
            {8'h00}, /* 0xd3d4 */
            {8'h00}, /* 0xd3d3 */
            {8'h00}, /* 0xd3d2 */
            {8'h00}, /* 0xd3d1 */
            {8'h00}, /* 0xd3d0 */
            {8'h00}, /* 0xd3cf */
            {8'h00}, /* 0xd3ce */
            {8'h00}, /* 0xd3cd */
            {8'h00}, /* 0xd3cc */
            {8'h00}, /* 0xd3cb */
            {8'h00}, /* 0xd3ca */
            {8'h00}, /* 0xd3c9 */
            {8'h00}, /* 0xd3c8 */
            {8'h00}, /* 0xd3c7 */
            {8'h00}, /* 0xd3c6 */
            {8'h00}, /* 0xd3c5 */
            {8'h00}, /* 0xd3c4 */
            {8'h00}, /* 0xd3c3 */
            {8'h00}, /* 0xd3c2 */
            {8'h00}, /* 0xd3c1 */
            {8'h00}, /* 0xd3c0 */
            {8'h00}, /* 0xd3bf */
            {8'h00}, /* 0xd3be */
            {8'h00}, /* 0xd3bd */
            {8'h00}, /* 0xd3bc */
            {8'h00}, /* 0xd3bb */
            {8'h00}, /* 0xd3ba */
            {8'h00}, /* 0xd3b9 */
            {8'h00}, /* 0xd3b8 */
            {8'h00}, /* 0xd3b7 */
            {8'h00}, /* 0xd3b6 */
            {8'h00}, /* 0xd3b5 */
            {8'h00}, /* 0xd3b4 */
            {8'h00}, /* 0xd3b3 */
            {8'h00}, /* 0xd3b2 */
            {8'h00}, /* 0xd3b1 */
            {8'h00}, /* 0xd3b0 */
            {8'h00}, /* 0xd3af */
            {8'h00}, /* 0xd3ae */
            {8'h00}, /* 0xd3ad */
            {8'h00}, /* 0xd3ac */
            {8'h00}, /* 0xd3ab */
            {8'h00}, /* 0xd3aa */
            {8'h00}, /* 0xd3a9 */
            {8'h00}, /* 0xd3a8 */
            {8'h00}, /* 0xd3a7 */
            {8'h00}, /* 0xd3a6 */
            {8'h00}, /* 0xd3a5 */
            {8'h00}, /* 0xd3a4 */
            {8'h00}, /* 0xd3a3 */
            {8'h00}, /* 0xd3a2 */
            {8'h00}, /* 0xd3a1 */
            {8'h00}, /* 0xd3a0 */
            {8'h00}, /* 0xd39f */
            {8'h00}, /* 0xd39e */
            {8'h00}, /* 0xd39d */
            {8'h00}, /* 0xd39c */
            {8'h00}, /* 0xd39b */
            {8'h00}, /* 0xd39a */
            {8'h00}, /* 0xd399 */
            {8'h00}, /* 0xd398 */
            {8'h00}, /* 0xd397 */
            {8'h00}, /* 0xd396 */
            {8'h00}, /* 0xd395 */
            {8'h00}, /* 0xd394 */
            {8'h00}, /* 0xd393 */
            {8'h00}, /* 0xd392 */
            {8'h00}, /* 0xd391 */
            {8'h00}, /* 0xd390 */
            {8'h00}, /* 0xd38f */
            {8'h00}, /* 0xd38e */
            {8'h00}, /* 0xd38d */
            {8'h00}, /* 0xd38c */
            {8'h00}, /* 0xd38b */
            {8'h00}, /* 0xd38a */
            {8'h00}, /* 0xd389 */
            {8'h00}, /* 0xd388 */
            {8'h00}, /* 0xd387 */
            {8'h00}, /* 0xd386 */
            {8'h00}, /* 0xd385 */
            {8'h00}, /* 0xd384 */
            {8'h00}, /* 0xd383 */
            {8'h00}, /* 0xd382 */
            {8'h00}, /* 0xd381 */
            {8'h00}, /* 0xd380 */
            {8'h00}, /* 0xd37f */
            {8'h00}, /* 0xd37e */
            {8'h00}, /* 0xd37d */
            {8'h00}, /* 0xd37c */
            {8'h00}, /* 0xd37b */
            {8'h00}, /* 0xd37a */
            {8'h00}, /* 0xd379 */
            {8'h00}, /* 0xd378 */
            {8'h00}, /* 0xd377 */
            {8'h00}, /* 0xd376 */
            {8'h00}, /* 0xd375 */
            {8'h00}, /* 0xd374 */
            {8'h00}, /* 0xd373 */
            {8'h00}, /* 0xd372 */
            {8'h00}, /* 0xd371 */
            {8'h00}, /* 0xd370 */
            {8'h00}, /* 0xd36f */
            {8'h00}, /* 0xd36e */
            {8'h00}, /* 0xd36d */
            {8'h00}, /* 0xd36c */
            {8'h00}, /* 0xd36b */
            {8'h00}, /* 0xd36a */
            {8'h00}, /* 0xd369 */
            {8'h00}, /* 0xd368 */
            {8'h00}, /* 0xd367 */
            {8'h00}, /* 0xd366 */
            {8'h00}, /* 0xd365 */
            {8'h00}, /* 0xd364 */
            {8'h00}, /* 0xd363 */
            {8'h00}, /* 0xd362 */
            {8'h00}, /* 0xd361 */
            {8'h00}, /* 0xd360 */
            {8'h00}, /* 0xd35f */
            {8'h00}, /* 0xd35e */
            {8'h00}, /* 0xd35d */
            {8'h00}, /* 0xd35c */
            {8'h00}, /* 0xd35b */
            {8'h00}, /* 0xd35a */
            {8'h00}, /* 0xd359 */
            {8'h00}, /* 0xd358 */
            {8'h00}, /* 0xd357 */
            {8'h00}, /* 0xd356 */
            {8'h00}, /* 0xd355 */
            {8'h00}, /* 0xd354 */
            {8'h00}, /* 0xd353 */
            {8'h00}, /* 0xd352 */
            {8'h00}, /* 0xd351 */
            {8'h00}, /* 0xd350 */
            {8'h00}, /* 0xd34f */
            {8'h00}, /* 0xd34e */
            {8'h00}, /* 0xd34d */
            {8'h00}, /* 0xd34c */
            {8'h00}, /* 0xd34b */
            {8'h00}, /* 0xd34a */
            {8'h00}, /* 0xd349 */
            {8'h00}, /* 0xd348 */
            {8'h00}, /* 0xd347 */
            {8'h00}, /* 0xd346 */
            {8'h00}, /* 0xd345 */
            {8'h00}, /* 0xd344 */
            {8'h00}, /* 0xd343 */
            {8'h00}, /* 0xd342 */
            {8'h00}, /* 0xd341 */
            {8'h00}, /* 0xd340 */
            {8'h00}, /* 0xd33f */
            {8'h00}, /* 0xd33e */
            {8'h00}, /* 0xd33d */
            {8'h00}, /* 0xd33c */
            {8'h00}, /* 0xd33b */
            {8'h00}, /* 0xd33a */
            {8'h00}, /* 0xd339 */
            {8'h00}, /* 0xd338 */
            {8'h00}, /* 0xd337 */
            {8'h00}, /* 0xd336 */
            {8'h00}, /* 0xd335 */
            {8'h00}, /* 0xd334 */
            {8'h00}, /* 0xd333 */
            {8'h00}, /* 0xd332 */
            {8'h00}, /* 0xd331 */
            {8'h00}, /* 0xd330 */
            {8'h00}, /* 0xd32f */
            {8'h00}, /* 0xd32e */
            {8'h00}, /* 0xd32d */
            {8'h00}, /* 0xd32c */
            {8'h00}, /* 0xd32b */
            {8'h00}, /* 0xd32a */
            {8'h00}, /* 0xd329 */
            {8'h00}, /* 0xd328 */
            {8'h00}, /* 0xd327 */
            {8'h00}, /* 0xd326 */
            {8'h00}, /* 0xd325 */
            {8'h00}, /* 0xd324 */
            {8'h00}, /* 0xd323 */
            {8'h00}, /* 0xd322 */
            {8'h00}, /* 0xd321 */
            {8'h00}, /* 0xd320 */
            {8'h00}, /* 0xd31f */
            {8'h00}, /* 0xd31e */
            {8'h00}, /* 0xd31d */
            {8'h00}, /* 0xd31c */
            {8'h00}, /* 0xd31b */
            {8'h00}, /* 0xd31a */
            {8'h00}, /* 0xd319 */
            {8'h00}, /* 0xd318 */
            {8'h00}, /* 0xd317 */
            {8'h00}, /* 0xd316 */
            {8'h00}, /* 0xd315 */
            {8'h00}, /* 0xd314 */
            {8'h00}, /* 0xd313 */
            {8'h00}, /* 0xd312 */
            {8'h00}, /* 0xd311 */
            {8'h00}, /* 0xd310 */
            {8'h00}, /* 0xd30f */
            {8'h00}, /* 0xd30e */
            {8'h00}, /* 0xd30d */
            {8'h00}, /* 0xd30c */
            {8'h00}, /* 0xd30b */
            {8'h00}, /* 0xd30a */
            {8'h00}, /* 0xd309 */
            {8'h00}, /* 0xd308 */
            {8'h00}, /* 0xd307 */
            {8'h00}, /* 0xd306 */
            {8'h00}, /* 0xd305 */
            {8'h00}, /* 0xd304 */
            {8'h00}, /* 0xd303 */
            {8'h00}, /* 0xd302 */
            {8'h00}, /* 0xd301 */
            {8'h00}, /* 0xd300 */
            {8'h00}, /* 0xd2ff */
            {8'h00}, /* 0xd2fe */
            {8'h00}, /* 0xd2fd */
            {8'h00}, /* 0xd2fc */
            {8'h00}, /* 0xd2fb */
            {8'h00}, /* 0xd2fa */
            {8'h00}, /* 0xd2f9 */
            {8'h00}, /* 0xd2f8 */
            {8'h00}, /* 0xd2f7 */
            {8'h00}, /* 0xd2f6 */
            {8'h00}, /* 0xd2f5 */
            {8'h00}, /* 0xd2f4 */
            {8'h00}, /* 0xd2f3 */
            {8'h00}, /* 0xd2f2 */
            {8'h00}, /* 0xd2f1 */
            {8'h00}, /* 0xd2f0 */
            {8'h00}, /* 0xd2ef */
            {8'h00}, /* 0xd2ee */
            {8'h00}, /* 0xd2ed */
            {8'h00}, /* 0xd2ec */
            {8'h00}, /* 0xd2eb */
            {8'h00}, /* 0xd2ea */
            {8'h00}, /* 0xd2e9 */
            {8'h00}, /* 0xd2e8 */
            {8'h00}, /* 0xd2e7 */
            {8'h00}, /* 0xd2e6 */
            {8'h00}, /* 0xd2e5 */
            {8'h00}, /* 0xd2e4 */
            {8'h00}, /* 0xd2e3 */
            {8'h00}, /* 0xd2e2 */
            {8'h00}, /* 0xd2e1 */
            {8'h00}, /* 0xd2e0 */
            {8'h00}, /* 0xd2df */
            {8'h00}, /* 0xd2de */
            {8'h00}, /* 0xd2dd */
            {8'h00}, /* 0xd2dc */
            {8'h00}, /* 0xd2db */
            {8'h00}, /* 0xd2da */
            {8'h00}, /* 0xd2d9 */
            {8'h00}, /* 0xd2d8 */
            {8'h00}, /* 0xd2d7 */
            {8'h00}, /* 0xd2d6 */
            {8'h00}, /* 0xd2d5 */
            {8'h00}, /* 0xd2d4 */
            {8'h00}, /* 0xd2d3 */
            {8'h00}, /* 0xd2d2 */
            {8'h00}, /* 0xd2d1 */
            {8'h00}, /* 0xd2d0 */
            {8'h00}, /* 0xd2cf */
            {8'h00}, /* 0xd2ce */
            {8'h00}, /* 0xd2cd */
            {8'h00}, /* 0xd2cc */
            {8'h00}, /* 0xd2cb */
            {8'h00}, /* 0xd2ca */
            {8'h00}, /* 0xd2c9 */
            {8'h00}, /* 0xd2c8 */
            {8'h00}, /* 0xd2c7 */
            {8'h00}, /* 0xd2c6 */
            {8'h00}, /* 0xd2c5 */
            {8'h00}, /* 0xd2c4 */
            {8'h00}, /* 0xd2c3 */
            {8'h00}, /* 0xd2c2 */
            {8'h00}, /* 0xd2c1 */
            {8'h00}, /* 0xd2c0 */
            {8'h00}, /* 0xd2bf */
            {8'h00}, /* 0xd2be */
            {8'h00}, /* 0xd2bd */
            {8'h00}, /* 0xd2bc */
            {8'h00}, /* 0xd2bb */
            {8'h00}, /* 0xd2ba */
            {8'h00}, /* 0xd2b9 */
            {8'h00}, /* 0xd2b8 */
            {8'h00}, /* 0xd2b7 */
            {8'h00}, /* 0xd2b6 */
            {8'h00}, /* 0xd2b5 */
            {8'h00}, /* 0xd2b4 */
            {8'h00}, /* 0xd2b3 */
            {8'h00}, /* 0xd2b2 */
            {8'h00}, /* 0xd2b1 */
            {8'h00}, /* 0xd2b0 */
            {8'h00}, /* 0xd2af */
            {8'h00}, /* 0xd2ae */
            {8'h00}, /* 0xd2ad */
            {8'h00}, /* 0xd2ac */
            {8'h00}, /* 0xd2ab */
            {8'h00}, /* 0xd2aa */
            {8'h00}, /* 0xd2a9 */
            {8'h00}, /* 0xd2a8 */
            {8'h00}, /* 0xd2a7 */
            {8'h00}, /* 0xd2a6 */
            {8'h00}, /* 0xd2a5 */
            {8'h00}, /* 0xd2a4 */
            {8'h00}, /* 0xd2a3 */
            {8'h00}, /* 0xd2a2 */
            {8'h00}, /* 0xd2a1 */
            {8'h00}, /* 0xd2a0 */
            {8'h00}, /* 0xd29f */
            {8'h00}, /* 0xd29e */
            {8'h00}, /* 0xd29d */
            {8'h00}, /* 0xd29c */
            {8'h00}, /* 0xd29b */
            {8'h00}, /* 0xd29a */
            {8'h00}, /* 0xd299 */
            {8'h00}, /* 0xd298 */
            {8'h00}, /* 0xd297 */
            {8'h00}, /* 0xd296 */
            {8'h00}, /* 0xd295 */
            {8'h00}, /* 0xd294 */
            {8'h00}, /* 0xd293 */
            {8'h00}, /* 0xd292 */
            {8'h00}, /* 0xd291 */
            {8'h00}, /* 0xd290 */
            {8'h00}, /* 0xd28f */
            {8'h00}, /* 0xd28e */
            {8'h00}, /* 0xd28d */
            {8'h00}, /* 0xd28c */
            {8'h00}, /* 0xd28b */
            {8'h00}, /* 0xd28a */
            {8'h00}, /* 0xd289 */
            {8'h00}, /* 0xd288 */
            {8'h00}, /* 0xd287 */
            {8'h00}, /* 0xd286 */
            {8'h00}, /* 0xd285 */
            {8'h00}, /* 0xd284 */
            {8'h00}, /* 0xd283 */
            {8'h00}, /* 0xd282 */
            {8'h00}, /* 0xd281 */
            {8'h00}, /* 0xd280 */
            {8'h00}, /* 0xd27f */
            {8'h00}, /* 0xd27e */
            {8'h00}, /* 0xd27d */
            {8'h00}, /* 0xd27c */
            {8'h00}, /* 0xd27b */
            {8'h00}, /* 0xd27a */
            {8'h00}, /* 0xd279 */
            {8'h00}, /* 0xd278 */
            {8'h00}, /* 0xd277 */
            {8'h00}, /* 0xd276 */
            {8'h00}, /* 0xd275 */
            {8'h00}, /* 0xd274 */
            {8'h00}, /* 0xd273 */
            {8'h00}, /* 0xd272 */
            {8'h00}, /* 0xd271 */
            {8'h00}, /* 0xd270 */
            {8'h00}, /* 0xd26f */
            {8'h00}, /* 0xd26e */
            {8'h00}, /* 0xd26d */
            {8'h00}, /* 0xd26c */
            {8'h00}, /* 0xd26b */
            {8'h00}, /* 0xd26a */
            {8'h00}, /* 0xd269 */
            {8'h00}, /* 0xd268 */
            {8'h00}, /* 0xd267 */
            {8'h00}, /* 0xd266 */
            {8'h00}, /* 0xd265 */
            {8'h00}, /* 0xd264 */
            {8'h00}, /* 0xd263 */
            {8'h00}, /* 0xd262 */
            {8'h00}, /* 0xd261 */
            {8'h00}, /* 0xd260 */
            {8'h00}, /* 0xd25f */
            {8'h00}, /* 0xd25e */
            {8'h00}, /* 0xd25d */
            {8'h00}, /* 0xd25c */
            {8'h00}, /* 0xd25b */
            {8'h00}, /* 0xd25a */
            {8'h00}, /* 0xd259 */
            {8'h00}, /* 0xd258 */
            {8'h00}, /* 0xd257 */
            {8'h00}, /* 0xd256 */
            {8'h00}, /* 0xd255 */
            {8'h00}, /* 0xd254 */
            {8'h00}, /* 0xd253 */
            {8'h00}, /* 0xd252 */
            {8'h00}, /* 0xd251 */
            {8'h00}, /* 0xd250 */
            {8'h00}, /* 0xd24f */
            {8'h00}, /* 0xd24e */
            {8'h00}, /* 0xd24d */
            {8'h00}, /* 0xd24c */
            {8'h00}, /* 0xd24b */
            {8'h00}, /* 0xd24a */
            {8'h00}, /* 0xd249 */
            {8'h00}, /* 0xd248 */
            {8'h00}, /* 0xd247 */
            {8'h00}, /* 0xd246 */
            {8'h00}, /* 0xd245 */
            {8'h00}, /* 0xd244 */
            {8'h00}, /* 0xd243 */
            {8'h00}, /* 0xd242 */
            {8'h00}, /* 0xd241 */
            {8'h00}, /* 0xd240 */
            {8'h00}, /* 0xd23f */
            {8'h00}, /* 0xd23e */
            {8'h00}, /* 0xd23d */
            {8'h00}, /* 0xd23c */
            {8'h00}, /* 0xd23b */
            {8'h00}, /* 0xd23a */
            {8'h00}, /* 0xd239 */
            {8'h00}, /* 0xd238 */
            {8'h00}, /* 0xd237 */
            {8'h00}, /* 0xd236 */
            {8'h00}, /* 0xd235 */
            {8'h00}, /* 0xd234 */
            {8'h00}, /* 0xd233 */
            {8'h00}, /* 0xd232 */
            {8'h00}, /* 0xd231 */
            {8'h00}, /* 0xd230 */
            {8'h00}, /* 0xd22f */
            {8'h00}, /* 0xd22e */
            {8'h00}, /* 0xd22d */
            {8'h00}, /* 0xd22c */
            {8'h00}, /* 0xd22b */
            {8'h00}, /* 0xd22a */
            {8'h00}, /* 0xd229 */
            {8'h00}, /* 0xd228 */
            {8'h00}, /* 0xd227 */
            {8'h00}, /* 0xd226 */
            {8'h00}, /* 0xd225 */
            {8'h00}, /* 0xd224 */
            {8'h00}, /* 0xd223 */
            {8'h00}, /* 0xd222 */
            {8'h00}, /* 0xd221 */
            {8'h00}, /* 0xd220 */
            {8'h00}, /* 0xd21f */
            {8'h00}, /* 0xd21e */
            {8'h00}, /* 0xd21d */
            {8'h00}, /* 0xd21c */
            {8'h00}, /* 0xd21b */
            {8'h00}, /* 0xd21a */
            {8'h00}, /* 0xd219 */
            {8'h00}, /* 0xd218 */
            {8'h00}, /* 0xd217 */
            {8'h00}, /* 0xd216 */
            {8'h00}, /* 0xd215 */
            {8'h00}, /* 0xd214 */
            {8'h00}, /* 0xd213 */
            {8'h00}, /* 0xd212 */
            {8'h00}, /* 0xd211 */
            {8'h00}, /* 0xd210 */
            {8'h00}, /* 0xd20f */
            {8'h00}, /* 0xd20e */
            {8'h00}, /* 0xd20d */
            {8'h00}, /* 0xd20c */
            {8'h00}, /* 0xd20b */
            {8'h00}, /* 0xd20a */
            {8'h00}, /* 0xd209 */
            {8'h00}, /* 0xd208 */
            {8'h00}, /* 0xd207 */
            {8'h00}, /* 0xd206 */
            {8'h00}, /* 0xd205 */
            {8'h00}, /* 0xd204 */
            {8'h00}, /* 0xd203 */
            {8'h00}, /* 0xd202 */
            {8'h00}, /* 0xd201 */
            {8'h00}, /* 0xd200 */
            {8'h00}, /* 0xd1ff */
            {8'h00}, /* 0xd1fe */
            {8'h00}, /* 0xd1fd */
            {8'h00}, /* 0xd1fc */
            {8'h00}, /* 0xd1fb */
            {8'h00}, /* 0xd1fa */
            {8'h00}, /* 0xd1f9 */
            {8'h00}, /* 0xd1f8 */
            {8'h00}, /* 0xd1f7 */
            {8'h00}, /* 0xd1f6 */
            {8'h00}, /* 0xd1f5 */
            {8'h00}, /* 0xd1f4 */
            {8'h00}, /* 0xd1f3 */
            {8'h00}, /* 0xd1f2 */
            {8'h00}, /* 0xd1f1 */
            {8'h00}, /* 0xd1f0 */
            {8'h00}, /* 0xd1ef */
            {8'h00}, /* 0xd1ee */
            {8'h00}, /* 0xd1ed */
            {8'h00}, /* 0xd1ec */
            {8'h00}, /* 0xd1eb */
            {8'h00}, /* 0xd1ea */
            {8'h00}, /* 0xd1e9 */
            {8'h00}, /* 0xd1e8 */
            {8'h00}, /* 0xd1e7 */
            {8'h00}, /* 0xd1e6 */
            {8'h00}, /* 0xd1e5 */
            {8'h00}, /* 0xd1e4 */
            {8'h00}, /* 0xd1e3 */
            {8'h00}, /* 0xd1e2 */
            {8'h00}, /* 0xd1e1 */
            {8'h00}, /* 0xd1e0 */
            {8'h00}, /* 0xd1df */
            {8'h00}, /* 0xd1de */
            {8'h00}, /* 0xd1dd */
            {8'h00}, /* 0xd1dc */
            {8'h00}, /* 0xd1db */
            {8'h00}, /* 0xd1da */
            {8'h00}, /* 0xd1d9 */
            {8'h00}, /* 0xd1d8 */
            {8'h00}, /* 0xd1d7 */
            {8'h00}, /* 0xd1d6 */
            {8'h00}, /* 0xd1d5 */
            {8'h00}, /* 0xd1d4 */
            {8'h00}, /* 0xd1d3 */
            {8'h00}, /* 0xd1d2 */
            {8'h00}, /* 0xd1d1 */
            {8'h00}, /* 0xd1d0 */
            {8'h00}, /* 0xd1cf */
            {8'h00}, /* 0xd1ce */
            {8'h00}, /* 0xd1cd */
            {8'h00}, /* 0xd1cc */
            {8'h00}, /* 0xd1cb */
            {8'h00}, /* 0xd1ca */
            {8'h00}, /* 0xd1c9 */
            {8'h00}, /* 0xd1c8 */
            {8'h00}, /* 0xd1c7 */
            {8'h00}, /* 0xd1c6 */
            {8'h00}, /* 0xd1c5 */
            {8'h00}, /* 0xd1c4 */
            {8'h00}, /* 0xd1c3 */
            {8'h00}, /* 0xd1c2 */
            {8'h00}, /* 0xd1c1 */
            {8'h00}, /* 0xd1c0 */
            {8'h00}, /* 0xd1bf */
            {8'h00}, /* 0xd1be */
            {8'h00}, /* 0xd1bd */
            {8'h00}, /* 0xd1bc */
            {8'h00}, /* 0xd1bb */
            {8'h00}, /* 0xd1ba */
            {8'h00}, /* 0xd1b9 */
            {8'h00}, /* 0xd1b8 */
            {8'h00}, /* 0xd1b7 */
            {8'h00}, /* 0xd1b6 */
            {8'h00}, /* 0xd1b5 */
            {8'h00}, /* 0xd1b4 */
            {8'h00}, /* 0xd1b3 */
            {8'h00}, /* 0xd1b2 */
            {8'h00}, /* 0xd1b1 */
            {8'h00}, /* 0xd1b0 */
            {8'h00}, /* 0xd1af */
            {8'h00}, /* 0xd1ae */
            {8'h00}, /* 0xd1ad */
            {8'h00}, /* 0xd1ac */
            {8'h00}, /* 0xd1ab */
            {8'h00}, /* 0xd1aa */
            {8'h00}, /* 0xd1a9 */
            {8'h00}, /* 0xd1a8 */
            {8'h00}, /* 0xd1a7 */
            {8'h00}, /* 0xd1a6 */
            {8'h00}, /* 0xd1a5 */
            {8'h00}, /* 0xd1a4 */
            {8'h00}, /* 0xd1a3 */
            {8'h00}, /* 0xd1a2 */
            {8'h00}, /* 0xd1a1 */
            {8'h00}, /* 0xd1a0 */
            {8'h00}, /* 0xd19f */
            {8'h00}, /* 0xd19e */
            {8'h00}, /* 0xd19d */
            {8'h00}, /* 0xd19c */
            {8'h00}, /* 0xd19b */
            {8'h00}, /* 0xd19a */
            {8'h00}, /* 0xd199 */
            {8'h00}, /* 0xd198 */
            {8'h00}, /* 0xd197 */
            {8'h00}, /* 0xd196 */
            {8'h00}, /* 0xd195 */
            {8'h00}, /* 0xd194 */
            {8'h00}, /* 0xd193 */
            {8'h00}, /* 0xd192 */
            {8'h00}, /* 0xd191 */
            {8'h00}, /* 0xd190 */
            {8'h00}, /* 0xd18f */
            {8'h00}, /* 0xd18e */
            {8'h00}, /* 0xd18d */
            {8'h00}, /* 0xd18c */
            {8'h00}, /* 0xd18b */
            {8'h00}, /* 0xd18a */
            {8'h00}, /* 0xd189 */
            {8'h00}, /* 0xd188 */
            {8'h00}, /* 0xd187 */
            {8'h00}, /* 0xd186 */
            {8'h00}, /* 0xd185 */
            {8'h00}, /* 0xd184 */
            {8'h00}, /* 0xd183 */
            {8'h00}, /* 0xd182 */
            {8'h00}, /* 0xd181 */
            {8'h00}, /* 0xd180 */
            {8'h00}, /* 0xd17f */
            {8'h00}, /* 0xd17e */
            {8'h00}, /* 0xd17d */
            {8'h00}, /* 0xd17c */
            {8'h00}, /* 0xd17b */
            {8'h00}, /* 0xd17a */
            {8'h00}, /* 0xd179 */
            {8'h00}, /* 0xd178 */
            {8'h00}, /* 0xd177 */
            {8'h00}, /* 0xd176 */
            {8'h00}, /* 0xd175 */
            {8'h00}, /* 0xd174 */
            {8'h00}, /* 0xd173 */
            {8'h00}, /* 0xd172 */
            {8'h00}, /* 0xd171 */
            {8'h00}, /* 0xd170 */
            {8'h00}, /* 0xd16f */
            {8'h00}, /* 0xd16e */
            {8'h00}, /* 0xd16d */
            {8'h00}, /* 0xd16c */
            {8'h00}, /* 0xd16b */
            {8'h00}, /* 0xd16a */
            {8'h00}, /* 0xd169 */
            {8'h00}, /* 0xd168 */
            {8'h00}, /* 0xd167 */
            {8'h00}, /* 0xd166 */
            {8'h00}, /* 0xd165 */
            {8'h00}, /* 0xd164 */
            {8'h00}, /* 0xd163 */
            {8'h00}, /* 0xd162 */
            {8'h00}, /* 0xd161 */
            {8'h00}, /* 0xd160 */
            {8'h00}, /* 0xd15f */
            {8'h00}, /* 0xd15e */
            {8'h00}, /* 0xd15d */
            {8'h00}, /* 0xd15c */
            {8'h00}, /* 0xd15b */
            {8'h00}, /* 0xd15a */
            {8'h00}, /* 0xd159 */
            {8'h00}, /* 0xd158 */
            {8'h00}, /* 0xd157 */
            {8'h00}, /* 0xd156 */
            {8'h00}, /* 0xd155 */
            {8'h00}, /* 0xd154 */
            {8'h00}, /* 0xd153 */
            {8'h00}, /* 0xd152 */
            {8'h00}, /* 0xd151 */
            {8'h00}, /* 0xd150 */
            {8'h00}, /* 0xd14f */
            {8'h00}, /* 0xd14e */
            {8'h00}, /* 0xd14d */
            {8'h00}, /* 0xd14c */
            {8'h00}, /* 0xd14b */
            {8'h00}, /* 0xd14a */
            {8'h00}, /* 0xd149 */
            {8'h00}, /* 0xd148 */
            {8'h00}, /* 0xd147 */
            {8'h00}, /* 0xd146 */
            {8'h00}, /* 0xd145 */
            {8'h00}, /* 0xd144 */
            {8'h00}, /* 0xd143 */
            {8'h00}, /* 0xd142 */
            {8'h00}, /* 0xd141 */
            {8'h00}, /* 0xd140 */
            {8'h00}, /* 0xd13f */
            {8'h00}, /* 0xd13e */
            {8'h00}, /* 0xd13d */
            {8'h00}, /* 0xd13c */
            {8'h00}, /* 0xd13b */
            {8'h00}, /* 0xd13a */
            {8'h00}, /* 0xd139 */
            {8'h00}, /* 0xd138 */
            {8'h00}, /* 0xd137 */
            {8'h00}, /* 0xd136 */
            {8'h00}, /* 0xd135 */
            {8'h00}, /* 0xd134 */
            {8'h00}, /* 0xd133 */
            {8'h00}, /* 0xd132 */
            {8'h00}, /* 0xd131 */
            {8'h00}, /* 0xd130 */
            {8'h00}, /* 0xd12f */
            {8'h00}, /* 0xd12e */
            {8'h00}, /* 0xd12d */
            {8'h00}, /* 0xd12c */
            {8'h00}, /* 0xd12b */
            {8'h00}, /* 0xd12a */
            {8'h00}, /* 0xd129 */
            {8'h00}, /* 0xd128 */
            {8'h00}, /* 0xd127 */
            {8'h00}, /* 0xd126 */
            {8'h00}, /* 0xd125 */
            {8'h00}, /* 0xd124 */
            {8'h00}, /* 0xd123 */
            {8'h00}, /* 0xd122 */
            {8'h00}, /* 0xd121 */
            {8'h00}, /* 0xd120 */
            {8'h00}, /* 0xd11f */
            {8'h00}, /* 0xd11e */
            {8'h00}, /* 0xd11d */
            {8'h00}, /* 0xd11c */
            {8'h00}, /* 0xd11b */
            {8'h00}, /* 0xd11a */
            {8'h00}, /* 0xd119 */
            {8'h00}, /* 0xd118 */
            {8'h00}, /* 0xd117 */
            {8'h00}, /* 0xd116 */
            {8'h00}, /* 0xd115 */
            {8'h00}, /* 0xd114 */
            {8'h00}, /* 0xd113 */
            {8'h00}, /* 0xd112 */
            {8'h00}, /* 0xd111 */
            {8'h00}, /* 0xd110 */
            {8'h00}, /* 0xd10f */
            {8'h00}, /* 0xd10e */
            {8'h00}, /* 0xd10d */
            {8'h00}, /* 0xd10c */
            {8'h00}, /* 0xd10b */
            {8'h00}, /* 0xd10a */
            {8'h00}, /* 0xd109 */
            {8'h00}, /* 0xd108 */
            {8'h00}, /* 0xd107 */
            {8'h00}, /* 0xd106 */
            {8'h00}, /* 0xd105 */
            {8'h00}, /* 0xd104 */
            {8'h00}, /* 0xd103 */
            {8'h00}, /* 0xd102 */
            {8'h00}, /* 0xd101 */
            {8'h00}, /* 0xd100 */
            {8'h00}, /* 0xd0ff */
            {8'h00}, /* 0xd0fe */
            {8'h00}, /* 0xd0fd */
            {8'h00}, /* 0xd0fc */
            {8'h00}, /* 0xd0fb */
            {8'h00}, /* 0xd0fa */
            {8'h00}, /* 0xd0f9 */
            {8'h00}, /* 0xd0f8 */
            {8'h00}, /* 0xd0f7 */
            {8'h00}, /* 0xd0f6 */
            {8'h00}, /* 0xd0f5 */
            {8'h00}, /* 0xd0f4 */
            {8'h00}, /* 0xd0f3 */
            {8'h00}, /* 0xd0f2 */
            {8'h00}, /* 0xd0f1 */
            {8'h00}, /* 0xd0f0 */
            {8'h00}, /* 0xd0ef */
            {8'h00}, /* 0xd0ee */
            {8'h00}, /* 0xd0ed */
            {8'h00}, /* 0xd0ec */
            {8'h00}, /* 0xd0eb */
            {8'h00}, /* 0xd0ea */
            {8'h00}, /* 0xd0e9 */
            {8'h00}, /* 0xd0e8 */
            {8'h00}, /* 0xd0e7 */
            {8'h00}, /* 0xd0e6 */
            {8'h00}, /* 0xd0e5 */
            {8'h00}, /* 0xd0e4 */
            {8'h00}, /* 0xd0e3 */
            {8'h00}, /* 0xd0e2 */
            {8'h00}, /* 0xd0e1 */
            {8'h00}, /* 0xd0e0 */
            {8'h00}, /* 0xd0df */
            {8'h00}, /* 0xd0de */
            {8'h00}, /* 0xd0dd */
            {8'h00}, /* 0xd0dc */
            {8'h00}, /* 0xd0db */
            {8'h00}, /* 0xd0da */
            {8'h00}, /* 0xd0d9 */
            {8'h00}, /* 0xd0d8 */
            {8'h00}, /* 0xd0d7 */
            {8'h00}, /* 0xd0d6 */
            {8'h00}, /* 0xd0d5 */
            {8'h00}, /* 0xd0d4 */
            {8'h00}, /* 0xd0d3 */
            {8'h00}, /* 0xd0d2 */
            {8'h00}, /* 0xd0d1 */
            {8'h00}, /* 0xd0d0 */
            {8'h00}, /* 0xd0cf */
            {8'h00}, /* 0xd0ce */
            {8'h00}, /* 0xd0cd */
            {8'h00}, /* 0xd0cc */
            {8'h00}, /* 0xd0cb */
            {8'h00}, /* 0xd0ca */
            {8'h00}, /* 0xd0c9 */
            {8'h00}, /* 0xd0c8 */
            {8'h00}, /* 0xd0c7 */
            {8'h00}, /* 0xd0c6 */
            {8'h00}, /* 0xd0c5 */
            {8'h00}, /* 0xd0c4 */
            {8'h00}, /* 0xd0c3 */
            {8'h00}, /* 0xd0c2 */
            {8'h00}, /* 0xd0c1 */
            {8'h00}, /* 0xd0c0 */
            {8'h00}, /* 0xd0bf */
            {8'h00}, /* 0xd0be */
            {8'h00}, /* 0xd0bd */
            {8'h00}, /* 0xd0bc */
            {8'h00}, /* 0xd0bb */
            {8'h00}, /* 0xd0ba */
            {8'h00}, /* 0xd0b9 */
            {8'h00}, /* 0xd0b8 */
            {8'h00}, /* 0xd0b7 */
            {8'h00}, /* 0xd0b6 */
            {8'h00}, /* 0xd0b5 */
            {8'h00}, /* 0xd0b4 */
            {8'h00}, /* 0xd0b3 */
            {8'h00}, /* 0xd0b2 */
            {8'h00}, /* 0xd0b1 */
            {8'h00}, /* 0xd0b0 */
            {8'h00}, /* 0xd0af */
            {8'h00}, /* 0xd0ae */
            {8'h00}, /* 0xd0ad */
            {8'h00}, /* 0xd0ac */
            {8'h00}, /* 0xd0ab */
            {8'h00}, /* 0xd0aa */
            {8'h00}, /* 0xd0a9 */
            {8'h00}, /* 0xd0a8 */
            {8'h00}, /* 0xd0a7 */
            {8'h00}, /* 0xd0a6 */
            {8'h00}, /* 0xd0a5 */
            {8'h00}, /* 0xd0a4 */
            {8'h00}, /* 0xd0a3 */
            {8'h00}, /* 0xd0a2 */
            {8'h00}, /* 0xd0a1 */
            {8'h00}, /* 0xd0a0 */
            {8'h00}, /* 0xd09f */
            {8'h00}, /* 0xd09e */
            {8'h00}, /* 0xd09d */
            {8'h00}, /* 0xd09c */
            {8'h00}, /* 0xd09b */
            {8'h00}, /* 0xd09a */
            {8'h00}, /* 0xd099 */
            {8'h00}, /* 0xd098 */
            {8'h00}, /* 0xd097 */
            {8'h00}, /* 0xd096 */
            {8'h00}, /* 0xd095 */
            {8'h00}, /* 0xd094 */
            {8'h00}, /* 0xd093 */
            {8'h00}, /* 0xd092 */
            {8'h00}, /* 0xd091 */
            {8'h00}, /* 0xd090 */
            {8'h00}, /* 0xd08f */
            {8'h00}, /* 0xd08e */
            {8'h00}, /* 0xd08d */
            {8'h00}, /* 0xd08c */
            {8'h00}, /* 0xd08b */
            {8'h00}, /* 0xd08a */
            {8'h00}, /* 0xd089 */
            {8'h00}, /* 0xd088 */
            {8'h00}, /* 0xd087 */
            {8'h00}, /* 0xd086 */
            {8'h00}, /* 0xd085 */
            {8'h00}, /* 0xd084 */
            {8'h00}, /* 0xd083 */
            {8'h00}, /* 0xd082 */
            {8'h00}, /* 0xd081 */
            {8'h00}, /* 0xd080 */
            {8'h00}, /* 0xd07f */
            {8'h00}, /* 0xd07e */
            {8'h00}, /* 0xd07d */
            {8'h00}, /* 0xd07c */
            {8'h00}, /* 0xd07b */
            {8'h00}, /* 0xd07a */
            {8'h00}, /* 0xd079 */
            {8'h00}, /* 0xd078 */
            {8'h00}, /* 0xd077 */
            {8'h00}, /* 0xd076 */
            {8'h00}, /* 0xd075 */
            {8'h00}, /* 0xd074 */
            {8'h00}, /* 0xd073 */
            {8'h00}, /* 0xd072 */
            {8'h00}, /* 0xd071 */
            {8'h00}, /* 0xd070 */
            {8'h00}, /* 0xd06f */
            {8'h00}, /* 0xd06e */
            {8'h00}, /* 0xd06d */
            {8'h00}, /* 0xd06c */
            {8'h00}, /* 0xd06b */
            {8'h00}, /* 0xd06a */
            {8'h00}, /* 0xd069 */
            {8'h00}, /* 0xd068 */
            {8'h00}, /* 0xd067 */
            {8'h00}, /* 0xd066 */
            {8'h00}, /* 0xd065 */
            {8'h00}, /* 0xd064 */
            {8'h00}, /* 0xd063 */
            {8'h00}, /* 0xd062 */
            {8'h00}, /* 0xd061 */
            {8'h00}, /* 0xd060 */
            {8'h00}, /* 0xd05f */
            {8'h00}, /* 0xd05e */
            {8'h00}, /* 0xd05d */
            {8'h00}, /* 0xd05c */
            {8'h00}, /* 0xd05b */
            {8'h00}, /* 0xd05a */
            {8'h00}, /* 0xd059 */
            {8'h00}, /* 0xd058 */
            {8'h00}, /* 0xd057 */
            {8'h00}, /* 0xd056 */
            {8'h00}, /* 0xd055 */
            {8'h00}, /* 0xd054 */
            {8'h00}, /* 0xd053 */
            {8'h00}, /* 0xd052 */
            {8'h00}, /* 0xd051 */
            {8'h00}, /* 0xd050 */
            {8'h00}, /* 0xd04f */
            {8'h00}, /* 0xd04e */
            {8'h00}, /* 0xd04d */
            {8'h00}, /* 0xd04c */
            {8'h00}, /* 0xd04b */
            {8'h00}, /* 0xd04a */
            {8'h00}, /* 0xd049 */
            {8'h00}, /* 0xd048 */
            {8'h00}, /* 0xd047 */
            {8'h00}, /* 0xd046 */
            {8'h00}, /* 0xd045 */
            {8'h00}, /* 0xd044 */
            {8'h00}, /* 0xd043 */
            {8'h00}, /* 0xd042 */
            {8'h00}, /* 0xd041 */
            {8'h00}, /* 0xd040 */
            {8'h00}, /* 0xd03f */
            {8'h00}, /* 0xd03e */
            {8'h00}, /* 0xd03d */
            {8'h00}, /* 0xd03c */
            {8'h00}, /* 0xd03b */
            {8'h00}, /* 0xd03a */
            {8'h00}, /* 0xd039 */
            {8'h00}, /* 0xd038 */
            {8'h00}, /* 0xd037 */
            {8'h00}, /* 0xd036 */
            {8'h00}, /* 0xd035 */
            {8'h00}, /* 0xd034 */
            {8'h00}, /* 0xd033 */
            {8'h00}, /* 0xd032 */
            {8'h00}, /* 0xd031 */
            {8'h00}, /* 0xd030 */
            {8'h00}, /* 0xd02f */
            {8'h00}, /* 0xd02e */
            {8'h00}, /* 0xd02d */
            {8'h00}, /* 0xd02c */
            {8'h00}, /* 0xd02b */
            {8'h00}, /* 0xd02a */
            {8'h00}, /* 0xd029 */
            {8'h00}, /* 0xd028 */
            {8'h00}, /* 0xd027 */
            {8'h00}, /* 0xd026 */
            {8'h00}, /* 0xd025 */
            {8'h00}, /* 0xd024 */
            {8'h00}, /* 0xd023 */
            {8'h00}, /* 0xd022 */
            {8'h00}, /* 0xd021 */
            {8'h00}, /* 0xd020 */
            {8'h00}, /* 0xd01f */
            {8'h00}, /* 0xd01e */
            {8'h00}, /* 0xd01d */
            {8'h00}, /* 0xd01c */
            {8'h00}, /* 0xd01b */
            {8'h00}, /* 0xd01a */
            {8'h00}, /* 0xd019 */
            {8'h00}, /* 0xd018 */
            {8'h00}, /* 0xd017 */
            {8'h00}, /* 0xd016 */
            {8'h00}, /* 0xd015 */
            {8'h00}, /* 0xd014 */
            {8'h00}, /* 0xd013 */
            {8'h00}, /* 0xd012 */
            {8'h00}, /* 0xd011 */
            {8'h00}, /* 0xd010 */
            {8'h00}, /* 0xd00f */
            {8'h00}, /* 0xd00e */
            {8'h00}, /* 0xd00d */
            {8'h00}, /* 0xd00c */
            {8'h00}, /* 0xd00b */
            {8'h00}, /* 0xd00a */
            {8'h00}, /* 0xd009 */
            {8'h00}, /* 0xd008 */
            {8'h00}, /* 0xd007 */
            {8'h00}, /* 0xd006 */
            {8'h00}, /* 0xd005 */
            {8'h00}, /* 0xd004 */
            {8'h00}, /* 0xd003 */
            {8'h00}, /* 0xd002 */
            {8'h00}, /* 0xd001 */
            {8'h00}, /* 0xd000 */
            {8'h00}, /* 0xcfff */
            {8'h00}, /* 0xcffe */
            {8'h00}, /* 0xcffd */
            {8'h00}, /* 0xcffc */
            {8'h00}, /* 0xcffb */
            {8'h00}, /* 0xcffa */
            {8'h00}, /* 0xcff9 */
            {8'h00}, /* 0xcff8 */
            {8'h00}, /* 0xcff7 */
            {8'h00}, /* 0xcff6 */
            {8'h00}, /* 0xcff5 */
            {8'h00}, /* 0xcff4 */
            {8'h00}, /* 0xcff3 */
            {8'h00}, /* 0xcff2 */
            {8'h00}, /* 0xcff1 */
            {8'h00}, /* 0xcff0 */
            {8'h00}, /* 0xcfef */
            {8'h00}, /* 0xcfee */
            {8'h00}, /* 0xcfed */
            {8'h00}, /* 0xcfec */
            {8'h00}, /* 0xcfeb */
            {8'h00}, /* 0xcfea */
            {8'h00}, /* 0xcfe9 */
            {8'h00}, /* 0xcfe8 */
            {8'h00}, /* 0xcfe7 */
            {8'h00}, /* 0xcfe6 */
            {8'h00}, /* 0xcfe5 */
            {8'h00}, /* 0xcfe4 */
            {8'h00}, /* 0xcfe3 */
            {8'h00}, /* 0xcfe2 */
            {8'h00}, /* 0xcfe1 */
            {8'h00}, /* 0xcfe0 */
            {8'h00}, /* 0xcfdf */
            {8'h00}, /* 0xcfde */
            {8'h00}, /* 0xcfdd */
            {8'h00}, /* 0xcfdc */
            {8'h00}, /* 0xcfdb */
            {8'h00}, /* 0xcfda */
            {8'h00}, /* 0xcfd9 */
            {8'h00}, /* 0xcfd8 */
            {8'h00}, /* 0xcfd7 */
            {8'h00}, /* 0xcfd6 */
            {8'h00}, /* 0xcfd5 */
            {8'h00}, /* 0xcfd4 */
            {8'h00}, /* 0xcfd3 */
            {8'h00}, /* 0xcfd2 */
            {8'h00}, /* 0xcfd1 */
            {8'h00}, /* 0xcfd0 */
            {8'h00}, /* 0xcfcf */
            {8'h00}, /* 0xcfce */
            {8'h00}, /* 0xcfcd */
            {8'h00}, /* 0xcfcc */
            {8'h00}, /* 0xcfcb */
            {8'h00}, /* 0xcfca */
            {8'h00}, /* 0xcfc9 */
            {8'h00}, /* 0xcfc8 */
            {8'h00}, /* 0xcfc7 */
            {8'h00}, /* 0xcfc6 */
            {8'h00}, /* 0xcfc5 */
            {8'h00}, /* 0xcfc4 */
            {8'h00}, /* 0xcfc3 */
            {8'h00}, /* 0xcfc2 */
            {8'h00}, /* 0xcfc1 */
            {8'h00}, /* 0xcfc0 */
            {8'h00}, /* 0xcfbf */
            {8'h00}, /* 0xcfbe */
            {8'h00}, /* 0xcfbd */
            {8'h00}, /* 0xcfbc */
            {8'h00}, /* 0xcfbb */
            {8'h00}, /* 0xcfba */
            {8'h00}, /* 0xcfb9 */
            {8'h00}, /* 0xcfb8 */
            {8'h00}, /* 0xcfb7 */
            {8'h00}, /* 0xcfb6 */
            {8'h00}, /* 0xcfb5 */
            {8'h00}, /* 0xcfb4 */
            {8'h00}, /* 0xcfb3 */
            {8'h00}, /* 0xcfb2 */
            {8'h00}, /* 0xcfb1 */
            {8'h00}, /* 0xcfb0 */
            {8'h00}, /* 0xcfaf */
            {8'h00}, /* 0xcfae */
            {8'h00}, /* 0xcfad */
            {8'h00}, /* 0xcfac */
            {8'h00}, /* 0xcfab */
            {8'h00}, /* 0xcfaa */
            {8'h00}, /* 0xcfa9 */
            {8'h00}, /* 0xcfa8 */
            {8'h00}, /* 0xcfa7 */
            {8'h00}, /* 0xcfa6 */
            {8'h00}, /* 0xcfa5 */
            {8'h00}, /* 0xcfa4 */
            {8'h00}, /* 0xcfa3 */
            {8'h00}, /* 0xcfa2 */
            {8'h00}, /* 0xcfa1 */
            {8'h00}, /* 0xcfa0 */
            {8'h00}, /* 0xcf9f */
            {8'h00}, /* 0xcf9e */
            {8'h00}, /* 0xcf9d */
            {8'h00}, /* 0xcf9c */
            {8'h00}, /* 0xcf9b */
            {8'h00}, /* 0xcf9a */
            {8'h00}, /* 0xcf99 */
            {8'h00}, /* 0xcf98 */
            {8'h00}, /* 0xcf97 */
            {8'h00}, /* 0xcf96 */
            {8'h00}, /* 0xcf95 */
            {8'h00}, /* 0xcf94 */
            {8'h00}, /* 0xcf93 */
            {8'h00}, /* 0xcf92 */
            {8'h00}, /* 0xcf91 */
            {8'h00}, /* 0xcf90 */
            {8'h00}, /* 0xcf8f */
            {8'h00}, /* 0xcf8e */
            {8'h00}, /* 0xcf8d */
            {8'h00}, /* 0xcf8c */
            {8'h00}, /* 0xcf8b */
            {8'h00}, /* 0xcf8a */
            {8'h00}, /* 0xcf89 */
            {8'h00}, /* 0xcf88 */
            {8'h00}, /* 0xcf87 */
            {8'h00}, /* 0xcf86 */
            {8'h00}, /* 0xcf85 */
            {8'h00}, /* 0xcf84 */
            {8'h00}, /* 0xcf83 */
            {8'h00}, /* 0xcf82 */
            {8'h00}, /* 0xcf81 */
            {8'h00}, /* 0xcf80 */
            {8'h00}, /* 0xcf7f */
            {8'h00}, /* 0xcf7e */
            {8'h00}, /* 0xcf7d */
            {8'h00}, /* 0xcf7c */
            {8'h00}, /* 0xcf7b */
            {8'h00}, /* 0xcf7a */
            {8'h00}, /* 0xcf79 */
            {8'h00}, /* 0xcf78 */
            {8'h00}, /* 0xcf77 */
            {8'h00}, /* 0xcf76 */
            {8'h00}, /* 0xcf75 */
            {8'h00}, /* 0xcf74 */
            {8'h00}, /* 0xcf73 */
            {8'h00}, /* 0xcf72 */
            {8'h00}, /* 0xcf71 */
            {8'h00}, /* 0xcf70 */
            {8'h00}, /* 0xcf6f */
            {8'h00}, /* 0xcf6e */
            {8'h00}, /* 0xcf6d */
            {8'h00}, /* 0xcf6c */
            {8'h00}, /* 0xcf6b */
            {8'h00}, /* 0xcf6a */
            {8'h00}, /* 0xcf69 */
            {8'h00}, /* 0xcf68 */
            {8'h00}, /* 0xcf67 */
            {8'h00}, /* 0xcf66 */
            {8'h00}, /* 0xcf65 */
            {8'h00}, /* 0xcf64 */
            {8'h00}, /* 0xcf63 */
            {8'h00}, /* 0xcf62 */
            {8'h00}, /* 0xcf61 */
            {8'h00}, /* 0xcf60 */
            {8'h00}, /* 0xcf5f */
            {8'h00}, /* 0xcf5e */
            {8'h00}, /* 0xcf5d */
            {8'h00}, /* 0xcf5c */
            {8'h00}, /* 0xcf5b */
            {8'h00}, /* 0xcf5a */
            {8'h00}, /* 0xcf59 */
            {8'h00}, /* 0xcf58 */
            {8'h00}, /* 0xcf57 */
            {8'h00}, /* 0xcf56 */
            {8'h00}, /* 0xcf55 */
            {8'h00}, /* 0xcf54 */
            {8'h00}, /* 0xcf53 */
            {8'h00}, /* 0xcf52 */
            {8'h00}, /* 0xcf51 */
            {8'h00}, /* 0xcf50 */
            {8'h00}, /* 0xcf4f */
            {8'h00}, /* 0xcf4e */
            {8'h00}, /* 0xcf4d */
            {8'h00}, /* 0xcf4c */
            {8'h00}, /* 0xcf4b */
            {8'h00}, /* 0xcf4a */
            {8'h00}, /* 0xcf49 */
            {8'h00}, /* 0xcf48 */
            {8'h00}, /* 0xcf47 */
            {8'h00}, /* 0xcf46 */
            {8'h00}, /* 0xcf45 */
            {8'h00}, /* 0xcf44 */
            {8'h00}, /* 0xcf43 */
            {8'h00}, /* 0xcf42 */
            {8'h00}, /* 0xcf41 */
            {8'h00}, /* 0xcf40 */
            {8'h00}, /* 0xcf3f */
            {8'h00}, /* 0xcf3e */
            {8'h00}, /* 0xcf3d */
            {8'h00}, /* 0xcf3c */
            {8'h00}, /* 0xcf3b */
            {8'h00}, /* 0xcf3a */
            {8'h00}, /* 0xcf39 */
            {8'h00}, /* 0xcf38 */
            {8'h00}, /* 0xcf37 */
            {8'h00}, /* 0xcf36 */
            {8'h00}, /* 0xcf35 */
            {8'h00}, /* 0xcf34 */
            {8'h00}, /* 0xcf33 */
            {8'h00}, /* 0xcf32 */
            {8'h00}, /* 0xcf31 */
            {8'h00}, /* 0xcf30 */
            {8'h00}, /* 0xcf2f */
            {8'h00}, /* 0xcf2e */
            {8'h00}, /* 0xcf2d */
            {8'h00}, /* 0xcf2c */
            {8'h00}, /* 0xcf2b */
            {8'h00}, /* 0xcf2a */
            {8'h00}, /* 0xcf29 */
            {8'h00}, /* 0xcf28 */
            {8'h00}, /* 0xcf27 */
            {8'h00}, /* 0xcf26 */
            {8'h00}, /* 0xcf25 */
            {8'h00}, /* 0xcf24 */
            {8'h00}, /* 0xcf23 */
            {8'h00}, /* 0xcf22 */
            {8'h00}, /* 0xcf21 */
            {8'h00}, /* 0xcf20 */
            {8'h00}, /* 0xcf1f */
            {8'h00}, /* 0xcf1e */
            {8'h00}, /* 0xcf1d */
            {8'h00}, /* 0xcf1c */
            {8'h00}, /* 0xcf1b */
            {8'h00}, /* 0xcf1a */
            {8'h00}, /* 0xcf19 */
            {8'h00}, /* 0xcf18 */
            {8'h00}, /* 0xcf17 */
            {8'h00}, /* 0xcf16 */
            {8'h00}, /* 0xcf15 */
            {8'h00}, /* 0xcf14 */
            {8'h00}, /* 0xcf13 */
            {8'h00}, /* 0xcf12 */
            {8'h00}, /* 0xcf11 */
            {8'h00}, /* 0xcf10 */
            {8'h00}, /* 0xcf0f */
            {8'h00}, /* 0xcf0e */
            {8'h00}, /* 0xcf0d */
            {8'h00}, /* 0xcf0c */
            {8'h00}, /* 0xcf0b */
            {8'h00}, /* 0xcf0a */
            {8'h00}, /* 0xcf09 */
            {8'h00}, /* 0xcf08 */
            {8'h00}, /* 0xcf07 */
            {8'h00}, /* 0xcf06 */
            {8'h00}, /* 0xcf05 */
            {8'h00}, /* 0xcf04 */
            {8'h00}, /* 0xcf03 */
            {8'h00}, /* 0xcf02 */
            {8'h00}, /* 0xcf01 */
            {8'h00}, /* 0xcf00 */
            {8'h00}, /* 0xceff */
            {8'h00}, /* 0xcefe */
            {8'h00}, /* 0xcefd */
            {8'h00}, /* 0xcefc */
            {8'h00}, /* 0xcefb */
            {8'h00}, /* 0xcefa */
            {8'h00}, /* 0xcef9 */
            {8'h00}, /* 0xcef8 */
            {8'h00}, /* 0xcef7 */
            {8'h00}, /* 0xcef6 */
            {8'h00}, /* 0xcef5 */
            {8'h00}, /* 0xcef4 */
            {8'h00}, /* 0xcef3 */
            {8'h00}, /* 0xcef2 */
            {8'h00}, /* 0xcef1 */
            {8'h00}, /* 0xcef0 */
            {8'h00}, /* 0xceef */
            {8'h00}, /* 0xceee */
            {8'h00}, /* 0xceed */
            {8'h00}, /* 0xceec */
            {8'h00}, /* 0xceeb */
            {8'h00}, /* 0xceea */
            {8'h00}, /* 0xcee9 */
            {8'h00}, /* 0xcee8 */
            {8'h00}, /* 0xcee7 */
            {8'h00}, /* 0xcee6 */
            {8'h00}, /* 0xcee5 */
            {8'h00}, /* 0xcee4 */
            {8'h00}, /* 0xcee3 */
            {8'h00}, /* 0xcee2 */
            {8'h00}, /* 0xcee1 */
            {8'h00}, /* 0xcee0 */
            {8'h00}, /* 0xcedf */
            {8'h00}, /* 0xcede */
            {8'h00}, /* 0xcedd */
            {8'h00}, /* 0xcedc */
            {8'h00}, /* 0xcedb */
            {8'h00}, /* 0xceda */
            {8'h00}, /* 0xced9 */
            {8'h00}, /* 0xced8 */
            {8'h00}, /* 0xced7 */
            {8'h00}, /* 0xced6 */
            {8'h00}, /* 0xced5 */
            {8'h00}, /* 0xced4 */
            {8'h00}, /* 0xced3 */
            {8'h00}, /* 0xced2 */
            {8'h00}, /* 0xced1 */
            {8'h00}, /* 0xced0 */
            {8'h00}, /* 0xcecf */
            {8'h00}, /* 0xcece */
            {8'h00}, /* 0xcecd */
            {8'h00}, /* 0xcecc */
            {8'h00}, /* 0xcecb */
            {8'h00}, /* 0xceca */
            {8'h00}, /* 0xcec9 */
            {8'h00}, /* 0xcec8 */
            {8'h00}, /* 0xcec7 */
            {8'h00}, /* 0xcec6 */
            {8'h00}, /* 0xcec5 */
            {8'h00}, /* 0xcec4 */
            {8'h00}, /* 0xcec3 */
            {8'h00}, /* 0xcec2 */
            {8'h00}, /* 0xcec1 */
            {8'h00}, /* 0xcec0 */
            {8'h00}, /* 0xcebf */
            {8'h00}, /* 0xcebe */
            {8'h00}, /* 0xcebd */
            {8'h00}, /* 0xcebc */
            {8'h00}, /* 0xcebb */
            {8'h00}, /* 0xceba */
            {8'h00}, /* 0xceb9 */
            {8'h00}, /* 0xceb8 */
            {8'h00}, /* 0xceb7 */
            {8'h00}, /* 0xceb6 */
            {8'h00}, /* 0xceb5 */
            {8'h00}, /* 0xceb4 */
            {8'h00}, /* 0xceb3 */
            {8'h00}, /* 0xceb2 */
            {8'h00}, /* 0xceb1 */
            {8'h00}, /* 0xceb0 */
            {8'h00}, /* 0xceaf */
            {8'h00}, /* 0xceae */
            {8'h00}, /* 0xcead */
            {8'h00}, /* 0xceac */
            {8'h00}, /* 0xceab */
            {8'h00}, /* 0xceaa */
            {8'h00}, /* 0xcea9 */
            {8'h00}, /* 0xcea8 */
            {8'h00}, /* 0xcea7 */
            {8'h00}, /* 0xcea6 */
            {8'h00}, /* 0xcea5 */
            {8'h00}, /* 0xcea4 */
            {8'h00}, /* 0xcea3 */
            {8'h00}, /* 0xcea2 */
            {8'h00}, /* 0xcea1 */
            {8'h00}, /* 0xcea0 */
            {8'h00}, /* 0xce9f */
            {8'h00}, /* 0xce9e */
            {8'h00}, /* 0xce9d */
            {8'h00}, /* 0xce9c */
            {8'h00}, /* 0xce9b */
            {8'h00}, /* 0xce9a */
            {8'h00}, /* 0xce99 */
            {8'h00}, /* 0xce98 */
            {8'h00}, /* 0xce97 */
            {8'h00}, /* 0xce96 */
            {8'h00}, /* 0xce95 */
            {8'h00}, /* 0xce94 */
            {8'h00}, /* 0xce93 */
            {8'h00}, /* 0xce92 */
            {8'h00}, /* 0xce91 */
            {8'h00}, /* 0xce90 */
            {8'h00}, /* 0xce8f */
            {8'h00}, /* 0xce8e */
            {8'h00}, /* 0xce8d */
            {8'h00}, /* 0xce8c */
            {8'h00}, /* 0xce8b */
            {8'h00}, /* 0xce8a */
            {8'h00}, /* 0xce89 */
            {8'h00}, /* 0xce88 */
            {8'h00}, /* 0xce87 */
            {8'h00}, /* 0xce86 */
            {8'h00}, /* 0xce85 */
            {8'h00}, /* 0xce84 */
            {8'h00}, /* 0xce83 */
            {8'h00}, /* 0xce82 */
            {8'h00}, /* 0xce81 */
            {8'h00}, /* 0xce80 */
            {8'h00}, /* 0xce7f */
            {8'h00}, /* 0xce7e */
            {8'h00}, /* 0xce7d */
            {8'h00}, /* 0xce7c */
            {8'h00}, /* 0xce7b */
            {8'h00}, /* 0xce7a */
            {8'h00}, /* 0xce79 */
            {8'h00}, /* 0xce78 */
            {8'h00}, /* 0xce77 */
            {8'h00}, /* 0xce76 */
            {8'h00}, /* 0xce75 */
            {8'h00}, /* 0xce74 */
            {8'h00}, /* 0xce73 */
            {8'h00}, /* 0xce72 */
            {8'h00}, /* 0xce71 */
            {8'h00}, /* 0xce70 */
            {8'h00}, /* 0xce6f */
            {8'h00}, /* 0xce6e */
            {8'h00}, /* 0xce6d */
            {8'h00}, /* 0xce6c */
            {8'h00}, /* 0xce6b */
            {8'h00}, /* 0xce6a */
            {8'h00}, /* 0xce69 */
            {8'h00}, /* 0xce68 */
            {8'h00}, /* 0xce67 */
            {8'h00}, /* 0xce66 */
            {8'h00}, /* 0xce65 */
            {8'h00}, /* 0xce64 */
            {8'h00}, /* 0xce63 */
            {8'h00}, /* 0xce62 */
            {8'h00}, /* 0xce61 */
            {8'h00}, /* 0xce60 */
            {8'h00}, /* 0xce5f */
            {8'h00}, /* 0xce5e */
            {8'h00}, /* 0xce5d */
            {8'h00}, /* 0xce5c */
            {8'h00}, /* 0xce5b */
            {8'h00}, /* 0xce5a */
            {8'h00}, /* 0xce59 */
            {8'h00}, /* 0xce58 */
            {8'h00}, /* 0xce57 */
            {8'h00}, /* 0xce56 */
            {8'h00}, /* 0xce55 */
            {8'h00}, /* 0xce54 */
            {8'h00}, /* 0xce53 */
            {8'h00}, /* 0xce52 */
            {8'h00}, /* 0xce51 */
            {8'h00}, /* 0xce50 */
            {8'h00}, /* 0xce4f */
            {8'h00}, /* 0xce4e */
            {8'h00}, /* 0xce4d */
            {8'h00}, /* 0xce4c */
            {8'h00}, /* 0xce4b */
            {8'h00}, /* 0xce4a */
            {8'h00}, /* 0xce49 */
            {8'h00}, /* 0xce48 */
            {8'h00}, /* 0xce47 */
            {8'h00}, /* 0xce46 */
            {8'h00}, /* 0xce45 */
            {8'h00}, /* 0xce44 */
            {8'h00}, /* 0xce43 */
            {8'h00}, /* 0xce42 */
            {8'h00}, /* 0xce41 */
            {8'h00}, /* 0xce40 */
            {8'h00}, /* 0xce3f */
            {8'h00}, /* 0xce3e */
            {8'h00}, /* 0xce3d */
            {8'h00}, /* 0xce3c */
            {8'h00}, /* 0xce3b */
            {8'h00}, /* 0xce3a */
            {8'h00}, /* 0xce39 */
            {8'h00}, /* 0xce38 */
            {8'h00}, /* 0xce37 */
            {8'h00}, /* 0xce36 */
            {8'h00}, /* 0xce35 */
            {8'h00}, /* 0xce34 */
            {8'h00}, /* 0xce33 */
            {8'h00}, /* 0xce32 */
            {8'h00}, /* 0xce31 */
            {8'h00}, /* 0xce30 */
            {8'h00}, /* 0xce2f */
            {8'h00}, /* 0xce2e */
            {8'h00}, /* 0xce2d */
            {8'h00}, /* 0xce2c */
            {8'h00}, /* 0xce2b */
            {8'h00}, /* 0xce2a */
            {8'h00}, /* 0xce29 */
            {8'h00}, /* 0xce28 */
            {8'h00}, /* 0xce27 */
            {8'h00}, /* 0xce26 */
            {8'h00}, /* 0xce25 */
            {8'h00}, /* 0xce24 */
            {8'h00}, /* 0xce23 */
            {8'h00}, /* 0xce22 */
            {8'h00}, /* 0xce21 */
            {8'h00}, /* 0xce20 */
            {8'h00}, /* 0xce1f */
            {8'h00}, /* 0xce1e */
            {8'h00}, /* 0xce1d */
            {8'h00}, /* 0xce1c */
            {8'h00}, /* 0xce1b */
            {8'h00}, /* 0xce1a */
            {8'h00}, /* 0xce19 */
            {8'h00}, /* 0xce18 */
            {8'h00}, /* 0xce17 */
            {8'h00}, /* 0xce16 */
            {8'h00}, /* 0xce15 */
            {8'h00}, /* 0xce14 */
            {8'h00}, /* 0xce13 */
            {8'h00}, /* 0xce12 */
            {8'h00}, /* 0xce11 */
            {8'h00}, /* 0xce10 */
            {8'h00}, /* 0xce0f */
            {8'h00}, /* 0xce0e */
            {8'h00}, /* 0xce0d */
            {8'h00}, /* 0xce0c */
            {8'h00}, /* 0xce0b */
            {8'h00}, /* 0xce0a */
            {8'h00}, /* 0xce09 */
            {8'h00}, /* 0xce08 */
            {8'h00}, /* 0xce07 */
            {8'h00}, /* 0xce06 */
            {8'h00}, /* 0xce05 */
            {8'h00}, /* 0xce04 */
            {8'h00}, /* 0xce03 */
            {8'h00}, /* 0xce02 */
            {8'h00}, /* 0xce01 */
            {8'h00}, /* 0xce00 */
            {8'h00}, /* 0xcdff */
            {8'h00}, /* 0xcdfe */
            {8'h00}, /* 0xcdfd */
            {8'h00}, /* 0xcdfc */
            {8'h00}, /* 0xcdfb */
            {8'h00}, /* 0xcdfa */
            {8'h00}, /* 0xcdf9 */
            {8'h00}, /* 0xcdf8 */
            {8'h00}, /* 0xcdf7 */
            {8'h00}, /* 0xcdf6 */
            {8'h00}, /* 0xcdf5 */
            {8'h00}, /* 0xcdf4 */
            {8'h00}, /* 0xcdf3 */
            {8'h00}, /* 0xcdf2 */
            {8'h00}, /* 0xcdf1 */
            {8'h00}, /* 0xcdf0 */
            {8'h00}, /* 0xcdef */
            {8'h00}, /* 0xcdee */
            {8'h00}, /* 0xcded */
            {8'h00}, /* 0xcdec */
            {8'h00}, /* 0xcdeb */
            {8'h00}, /* 0xcdea */
            {8'h00}, /* 0xcde9 */
            {8'h00}, /* 0xcde8 */
            {8'h00}, /* 0xcde7 */
            {8'h00}, /* 0xcde6 */
            {8'h00}, /* 0xcde5 */
            {8'h00}, /* 0xcde4 */
            {8'h00}, /* 0xcde3 */
            {8'h00}, /* 0xcde2 */
            {8'h00}, /* 0xcde1 */
            {8'h00}, /* 0xcde0 */
            {8'h00}, /* 0xcddf */
            {8'h00}, /* 0xcdde */
            {8'h00}, /* 0xcddd */
            {8'h00}, /* 0xcddc */
            {8'h00}, /* 0xcddb */
            {8'h00}, /* 0xcdda */
            {8'h00}, /* 0xcdd9 */
            {8'h00}, /* 0xcdd8 */
            {8'h00}, /* 0xcdd7 */
            {8'h00}, /* 0xcdd6 */
            {8'h00}, /* 0xcdd5 */
            {8'h00}, /* 0xcdd4 */
            {8'h00}, /* 0xcdd3 */
            {8'h00}, /* 0xcdd2 */
            {8'h00}, /* 0xcdd1 */
            {8'h00}, /* 0xcdd0 */
            {8'h00}, /* 0xcdcf */
            {8'h00}, /* 0xcdce */
            {8'h00}, /* 0xcdcd */
            {8'h00}, /* 0xcdcc */
            {8'h00}, /* 0xcdcb */
            {8'h00}, /* 0xcdca */
            {8'h00}, /* 0xcdc9 */
            {8'h00}, /* 0xcdc8 */
            {8'h00}, /* 0xcdc7 */
            {8'h00}, /* 0xcdc6 */
            {8'h00}, /* 0xcdc5 */
            {8'h00}, /* 0xcdc4 */
            {8'h00}, /* 0xcdc3 */
            {8'h00}, /* 0xcdc2 */
            {8'h00}, /* 0xcdc1 */
            {8'h00}, /* 0xcdc0 */
            {8'h00}, /* 0xcdbf */
            {8'h00}, /* 0xcdbe */
            {8'h00}, /* 0xcdbd */
            {8'h00}, /* 0xcdbc */
            {8'h00}, /* 0xcdbb */
            {8'h00}, /* 0xcdba */
            {8'h00}, /* 0xcdb9 */
            {8'h00}, /* 0xcdb8 */
            {8'h00}, /* 0xcdb7 */
            {8'h00}, /* 0xcdb6 */
            {8'h00}, /* 0xcdb5 */
            {8'h00}, /* 0xcdb4 */
            {8'h00}, /* 0xcdb3 */
            {8'h00}, /* 0xcdb2 */
            {8'h00}, /* 0xcdb1 */
            {8'h00}, /* 0xcdb0 */
            {8'h00}, /* 0xcdaf */
            {8'h00}, /* 0xcdae */
            {8'h00}, /* 0xcdad */
            {8'h00}, /* 0xcdac */
            {8'h00}, /* 0xcdab */
            {8'h00}, /* 0xcdaa */
            {8'h00}, /* 0xcda9 */
            {8'h00}, /* 0xcda8 */
            {8'h00}, /* 0xcda7 */
            {8'h00}, /* 0xcda6 */
            {8'h00}, /* 0xcda5 */
            {8'h00}, /* 0xcda4 */
            {8'h00}, /* 0xcda3 */
            {8'h00}, /* 0xcda2 */
            {8'h00}, /* 0xcda1 */
            {8'h00}, /* 0xcda0 */
            {8'h00}, /* 0xcd9f */
            {8'h00}, /* 0xcd9e */
            {8'h00}, /* 0xcd9d */
            {8'h00}, /* 0xcd9c */
            {8'h00}, /* 0xcd9b */
            {8'h00}, /* 0xcd9a */
            {8'h00}, /* 0xcd99 */
            {8'h00}, /* 0xcd98 */
            {8'h00}, /* 0xcd97 */
            {8'h00}, /* 0xcd96 */
            {8'h00}, /* 0xcd95 */
            {8'h00}, /* 0xcd94 */
            {8'h00}, /* 0xcd93 */
            {8'h00}, /* 0xcd92 */
            {8'h00}, /* 0xcd91 */
            {8'h00}, /* 0xcd90 */
            {8'h00}, /* 0xcd8f */
            {8'h00}, /* 0xcd8e */
            {8'h00}, /* 0xcd8d */
            {8'h00}, /* 0xcd8c */
            {8'h00}, /* 0xcd8b */
            {8'h00}, /* 0xcd8a */
            {8'h00}, /* 0xcd89 */
            {8'h00}, /* 0xcd88 */
            {8'h00}, /* 0xcd87 */
            {8'h00}, /* 0xcd86 */
            {8'h00}, /* 0xcd85 */
            {8'h00}, /* 0xcd84 */
            {8'h00}, /* 0xcd83 */
            {8'h00}, /* 0xcd82 */
            {8'h00}, /* 0xcd81 */
            {8'h00}, /* 0xcd80 */
            {8'h00}, /* 0xcd7f */
            {8'h00}, /* 0xcd7e */
            {8'h00}, /* 0xcd7d */
            {8'h00}, /* 0xcd7c */
            {8'h00}, /* 0xcd7b */
            {8'h00}, /* 0xcd7a */
            {8'h00}, /* 0xcd79 */
            {8'h00}, /* 0xcd78 */
            {8'h00}, /* 0xcd77 */
            {8'h00}, /* 0xcd76 */
            {8'h00}, /* 0xcd75 */
            {8'h00}, /* 0xcd74 */
            {8'h00}, /* 0xcd73 */
            {8'h00}, /* 0xcd72 */
            {8'h00}, /* 0xcd71 */
            {8'h00}, /* 0xcd70 */
            {8'h00}, /* 0xcd6f */
            {8'h00}, /* 0xcd6e */
            {8'h00}, /* 0xcd6d */
            {8'h00}, /* 0xcd6c */
            {8'h00}, /* 0xcd6b */
            {8'h00}, /* 0xcd6a */
            {8'h00}, /* 0xcd69 */
            {8'h00}, /* 0xcd68 */
            {8'h00}, /* 0xcd67 */
            {8'h00}, /* 0xcd66 */
            {8'h00}, /* 0xcd65 */
            {8'h00}, /* 0xcd64 */
            {8'h00}, /* 0xcd63 */
            {8'h00}, /* 0xcd62 */
            {8'h00}, /* 0xcd61 */
            {8'h00}, /* 0xcd60 */
            {8'h00}, /* 0xcd5f */
            {8'h00}, /* 0xcd5e */
            {8'h00}, /* 0xcd5d */
            {8'h00}, /* 0xcd5c */
            {8'h00}, /* 0xcd5b */
            {8'h00}, /* 0xcd5a */
            {8'h00}, /* 0xcd59 */
            {8'h00}, /* 0xcd58 */
            {8'h00}, /* 0xcd57 */
            {8'h00}, /* 0xcd56 */
            {8'h00}, /* 0xcd55 */
            {8'h00}, /* 0xcd54 */
            {8'h00}, /* 0xcd53 */
            {8'h00}, /* 0xcd52 */
            {8'h00}, /* 0xcd51 */
            {8'h00}, /* 0xcd50 */
            {8'h00}, /* 0xcd4f */
            {8'h00}, /* 0xcd4e */
            {8'h00}, /* 0xcd4d */
            {8'h00}, /* 0xcd4c */
            {8'h00}, /* 0xcd4b */
            {8'h00}, /* 0xcd4a */
            {8'h00}, /* 0xcd49 */
            {8'h00}, /* 0xcd48 */
            {8'h00}, /* 0xcd47 */
            {8'h00}, /* 0xcd46 */
            {8'h00}, /* 0xcd45 */
            {8'h00}, /* 0xcd44 */
            {8'h00}, /* 0xcd43 */
            {8'h00}, /* 0xcd42 */
            {8'h00}, /* 0xcd41 */
            {8'h00}, /* 0xcd40 */
            {8'h00}, /* 0xcd3f */
            {8'h00}, /* 0xcd3e */
            {8'h00}, /* 0xcd3d */
            {8'h00}, /* 0xcd3c */
            {8'h00}, /* 0xcd3b */
            {8'h00}, /* 0xcd3a */
            {8'h00}, /* 0xcd39 */
            {8'h00}, /* 0xcd38 */
            {8'h00}, /* 0xcd37 */
            {8'h00}, /* 0xcd36 */
            {8'h00}, /* 0xcd35 */
            {8'h00}, /* 0xcd34 */
            {8'h00}, /* 0xcd33 */
            {8'h00}, /* 0xcd32 */
            {8'h00}, /* 0xcd31 */
            {8'h00}, /* 0xcd30 */
            {8'h00}, /* 0xcd2f */
            {8'h00}, /* 0xcd2e */
            {8'h00}, /* 0xcd2d */
            {8'h00}, /* 0xcd2c */
            {8'h00}, /* 0xcd2b */
            {8'h00}, /* 0xcd2a */
            {8'h00}, /* 0xcd29 */
            {8'h00}, /* 0xcd28 */
            {8'h00}, /* 0xcd27 */
            {8'h00}, /* 0xcd26 */
            {8'h00}, /* 0xcd25 */
            {8'h00}, /* 0xcd24 */
            {8'h00}, /* 0xcd23 */
            {8'h00}, /* 0xcd22 */
            {8'h00}, /* 0xcd21 */
            {8'h00}, /* 0xcd20 */
            {8'h00}, /* 0xcd1f */
            {8'h00}, /* 0xcd1e */
            {8'h00}, /* 0xcd1d */
            {8'h00}, /* 0xcd1c */
            {8'h00}, /* 0xcd1b */
            {8'h00}, /* 0xcd1a */
            {8'h00}, /* 0xcd19 */
            {8'h00}, /* 0xcd18 */
            {8'h00}, /* 0xcd17 */
            {8'h00}, /* 0xcd16 */
            {8'h00}, /* 0xcd15 */
            {8'h00}, /* 0xcd14 */
            {8'h00}, /* 0xcd13 */
            {8'h00}, /* 0xcd12 */
            {8'h00}, /* 0xcd11 */
            {8'h00}, /* 0xcd10 */
            {8'h00}, /* 0xcd0f */
            {8'h00}, /* 0xcd0e */
            {8'h00}, /* 0xcd0d */
            {8'h00}, /* 0xcd0c */
            {8'h00}, /* 0xcd0b */
            {8'h00}, /* 0xcd0a */
            {8'h00}, /* 0xcd09 */
            {8'h00}, /* 0xcd08 */
            {8'h00}, /* 0xcd07 */
            {8'h00}, /* 0xcd06 */
            {8'h00}, /* 0xcd05 */
            {8'h00}, /* 0xcd04 */
            {8'h00}, /* 0xcd03 */
            {8'h00}, /* 0xcd02 */
            {8'h00}, /* 0xcd01 */
            {8'h00}, /* 0xcd00 */
            {8'h00}, /* 0xccff */
            {8'h00}, /* 0xccfe */
            {8'h00}, /* 0xccfd */
            {8'h00}, /* 0xccfc */
            {8'h00}, /* 0xccfb */
            {8'h00}, /* 0xccfa */
            {8'h00}, /* 0xccf9 */
            {8'h00}, /* 0xccf8 */
            {8'h00}, /* 0xccf7 */
            {8'h00}, /* 0xccf6 */
            {8'h00}, /* 0xccf5 */
            {8'h00}, /* 0xccf4 */
            {8'h00}, /* 0xccf3 */
            {8'h00}, /* 0xccf2 */
            {8'h00}, /* 0xccf1 */
            {8'h00}, /* 0xccf0 */
            {8'h00}, /* 0xccef */
            {8'h00}, /* 0xccee */
            {8'h00}, /* 0xcced */
            {8'h00}, /* 0xccec */
            {8'h00}, /* 0xcceb */
            {8'h00}, /* 0xccea */
            {8'h00}, /* 0xcce9 */
            {8'h00}, /* 0xcce8 */
            {8'h00}, /* 0xcce7 */
            {8'h00}, /* 0xcce6 */
            {8'h00}, /* 0xcce5 */
            {8'h00}, /* 0xcce4 */
            {8'h00}, /* 0xcce3 */
            {8'h00}, /* 0xcce2 */
            {8'h00}, /* 0xcce1 */
            {8'h00}, /* 0xcce0 */
            {8'h00}, /* 0xccdf */
            {8'h00}, /* 0xccde */
            {8'h00}, /* 0xccdd */
            {8'h00}, /* 0xccdc */
            {8'h00}, /* 0xccdb */
            {8'h00}, /* 0xccda */
            {8'h00}, /* 0xccd9 */
            {8'h00}, /* 0xccd8 */
            {8'h00}, /* 0xccd7 */
            {8'h00}, /* 0xccd6 */
            {8'h00}, /* 0xccd5 */
            {8'h00}, /* 0xccd4 */
            {8'h00}, /* 0xccd3 */
            {8'h00}, /* 0xccd2 */
            {8'h00}, /* 0xccd1 */
            {8'h00}, /* 0xccd0 */
            {8'h00}, /* 0xcccf */
            {8'h00}, /* 0xccce */
            {8'h00}, /* 0xcccd */
            {8'h00}, /* 0xcccc */
            {8'h00}, /* 0xcccb */
            {8'h00}, /* 0xccca */
            {8'h00}, /* 0xccc9 */
            {8'h00}, /* 0xccc8 */
            {8'h00}, /* 0xccc7 */
            {8'h00}, /* 0xccc6 */
            {8'h00}, /* 0xccc5 */
            {8'h00}, /* 0xccc4 */
            {8'h00}, /* 0xccc3 */
            {8'h00}, /* 0xccc2 */
            {8'h00}, /* 0xccc1 */
            {8'h00}, /* 0xccc0 */
            {8'h00}, /* 0xccbf */
            {8'h00}, /* 0xccbe */
            {8'h00}, /* 0xccbd */
            {8'h00}, /* 0xccbc */
            {8'h00}, /* 0xccbb */
            {8'h00}, /* 0xccba */
            {8'h00}, /* 0xccb9 */
            {8'h00}, /* 0xccb8 */
            {8'h00}, /* 0xccb7 */
            {8'h00}, /* 0xccb6 */
            {8'h00}, /* 0xccb5 */
            {8'h00}, /* 0xccb4 */
            {8'h00}, /* 0xccb3 */
            {8'h00}, /* 0xccb2 */
            {8'h00}, /* 0xccb1 */
            {8'h00}, /* 0xccb0 */
            {8'h00}, /* 0xccaf */
            {8'h00}, /* 0xccae */
            {8'h00}, /* 0xccad */
            {8'h00}, /* 0xccac */
            {8'h00}, /* 0xccab */
            {8'h00}, /* 0xccaa */
            {8'h00}, /* 0xcca9 */
            {8'h00}, /* 0xcca8 */
            {8'h00}, /* 0xcca7 */
            {8'h00}, /* 0xcca6 */
            {8'h00}, /* 0xcca5 */
            {8'h00}, /* 0xcca4 */
            {8'h00}, /* 0xcca3 */
            {8'h00}, /* 0xcca2 */
            {8'h00}, /* 0xcca1 */
            {8'h00}, /* 0xcca0 */
            {8'h00}, /* 0xcc9f */
            {8'h00}, /* 0xcc9e */
            {8'h00}, /* 0xcc9d */
            {8'h00}, /* 0xcc9c */
            {8'h00}, /* 0xcc9b */
            {8'h00}, /* 0xcc9a */
            {8'h00}, /* 0xcc99 */
            {8'h00}, /* 0xcc98 */
            {8'h00}, /* 0xcc97 */
            {8'h00}, /* 0xcc96 */
            {8'h00}, /* 0xcc95 */
            {8'h00}, /* 0xcc94 */
            {8'h00}, /* 0xcc93 */
            {8'h00}, /* 0xcc92 */
            {8'h00}, /* 0xcc91 */
            {8'h00}, /* 0xcc90 */
            {8'h00}, /* 0xcc8f */
            {8'h00}, /* 0xcc8e */
            {8'h00}, /* 0xcc8d */
            {8'h00}, /* 0xcc8c */
            {8'h00}, /* 0xcc8b */
            {8'h00}, /* 0xcc8a */
            {8'h00}, /* 0xcc89 */
            {8'h00}, /* 0xcc88 */
            {8'h00}, /* 0xcc87 */
            {8'h00}, /* 0xcc86 */
            {8'h00}, /* 0xcc85 */
            {8'h00}, /* 0xcc84 */
            {8'h00}, /* 0xcc83 */
            {8'h00}, /* 0xcc82 */
            {8'h00}, /* 0xcc81 */
            {8'h00}, /* 0xcc80 */
            {8'h00}, /* 0xcc7f */
            {8'h00}, /* 0xcc7e */
            {8'h00}, /* 0xcc7d */
            {8'h00}, /* 0xcc7c */
            {8'h00}, /* 0xcc7b */
            {8'h00}, /* 0xcc7a */
            {8'h00}, /* 0xcc79 */
            {8'h00}, /* 0xcc78 */
            {8'h00}, /* 0xcc77 */
            {8'h00}, /* 0xcc76 */
            {8'h00}, /* 0xcc75 */
            {8'h00}, /* 0xcc74 */
            {8'h00}, /* 0xcc73 */
            {8'h00}, /* 0xcc72 */
            {8'h00}, /* 0xcc71 */
            {8'h00}, /* 0xcc70 */
            {8'h00}, /* 0xcc6f */
            {8'h00}, /* 0xcc6e */
            {8'h00}, /* 0xcc6d */
            {8'h00}, /* 0xcc6c */
            {8'h00}, /* 0xcc6b */
            {8'h00}, /* 0xcc6a */
            {8'h00}, /* 0xcc69 */
            {8'h00}, /* 0xcc68 */
            {8'h00}, /* 0xcc67 */
            {8'h00}, /* 0xcc66 */
            {8'h00}, /* 0xcc65 */
            {8'h00}, /* 0xcc64 */
            {8'h00}, /* 0xcc63 */
            {8'h00}, /* 0xcc62 */
            {8'h00}, /* 0xcc61 */
            {8'h00}, /* 0xcc60 */
            {8'h00}, /* 0xcc5f */
            {8'h00}, /* 0xcc5e */
            {8'h00}, /* 0xcc5d */
            {8'h00}, /* 0xcc5c */
            {8'h00}, /* 0xcc5b */
            {8'h00}, /* 0xcc5a */
            {8'h00}, /* 0xcc59 */
            {8'h00}, /* 0xcc58 */
            {8'h00}, /* 0xcc57 */
            {8'h00}, /* 0xcc56 */
            {8'h00}, /* 0xcc55 */
            {8'h00}, /* 0xcc54 */
            {8'h00}, /* 0xcc53 */
            {8'h00}, /* 0xcc52 */
            {8'h00}, /* 0xcc51 */
            {8'h00}, /* 0xcc50 */
            {8'h00}, /* 0xcc4f */
            {8'h00}, /* 0xcc4e */
            {8'h00}, /* 0xcc4d */
            {8'h00}, /* 0xcc4c */
            {8'h00}, /* 0xcc4b */
            {8'h00}, /* 0xcc4a */
            {8'h00}, /* 0xcc49 */
            {8'h00}, /* 0xcc48 */
            {8'h00}, /* 0xcc47 */
            {8'h00}, /* 0xcc46 */
            {8'h00}, /* 0xcc45 */
            {8'h00}, /* 0xcc44 */
            {8'h00}, /* 0xcc43 */
            {8'h00}, /* 0xcc42 */
            {8'h00}, /* 0xcc41 */
            {8'h00}, /* 0xcc40 */
            {8'h00}, /* 0xcc3f */
            {8'h00}, /* 0xcc3e */
            {8'h00}, /* 0xcc3d */
            {8'h00}, /* 0xcc3c */
            {8'h00}, /* 0xcc3b */
            {8'h00}, /* 0xcc3a */
            {8'h00}, /* 0xcc39 */
            {8'h00}, /* 0xcc38 */
            {8'h00}, /* 0xcc37 */
            {8'h00}, /* 0xcc36 */
            {8'h00}, /* 0xcc35 */
            {8'h00}, /* 0xcc34 */
            {8'h00}, /* 0xcc33 */
            {8'h00}, /* 0xcc32 */
            {8'h00}, /* 0xcc31 */
            {8'h00}, /* 0xcc30 */
            {8'h00}, /* 0xcc2f */
            {8'h00}, /* 0xcc2e */
            {8'h00}, /* 0xcc2d */
            {8'h00}, /* 0xcc2c */
            {8'h00}, /* 0xcc2b */
            {8'h00}, /* 0xcc2a */
            {8'h00}, /* 0xcc29 */
            {8'h00}, /* 0xcc28 */
            {8'h00}, /* 0xcc27 */
            {8'h00}, /* 0xcc26 */
            {8'h00}, /* 0xcc25 */
            {8'h00}, /* 0xcc24 */
            {8'h00}, /* 0xcc23 */
            {8'h00}, /* 0xcc22 */
            {8'h00}, /* 0xcc21 */
            {8'h00}, /* 0xcc20 */
            {8'h00}, /* 0xcc1f */
            {8'h00}, /* 0xcc1e */
            {8'h00}, /* 0xcc1d */
            {8'h00}, /* 0xcc1c */
            {8'h00}, /* 0xcc1b */
            {8'h00}, /* 0xcc1a */
            {8'h00}, /* 0xcc19 */
            {8'h00}, /* 0xcc18 */
            {8'h00}, /* 0xcc17 */
            {8'h00}, /* 0xcc16 */
            {8'h00}, /* 0xcc15 */
            {8'h00}, /* 0xcc14 */
            {8'h00}, /* 0xcc13 */
            {8'h00}, /* 0xcc12 */
            {8'h00}, /* 0xcc11 */
            {8'h00}, /* 0xcc10 */
            {8'h00}, /* 0xcc0f */
            {8'h00}, /* 0xcc0e */
            {8'h00}, /* 0xcc0d */
            {8'h00}, /* 0xcc0c */
            {8'h00}, /* 0xcc0b */
            {8'h00}, /* 0xcc0a */
            {8'h00}, /* 0xcc09 */
            {8'h00}, /* 0xcc08 */
            {8'h00}, /* 0xcc07 */
            {8'h00}, /* 0xcc06 */
            {8'h00}, /* 0xcc05 */
            {8'h00}, /* 0xcc04 */
            {8'h00}, /* 0xcc03 */
            {8'h00}, /* 0xcc02 */
            {8'h00}, /* 0xcc01 */
            {8'h00}, /* 0xcc00 */
            {8'h00}, /* 0xcbff */
            {8'h00}, /* 0xcbfe */
            {8'h00}, /* 0xcbfd */
            {8'h00}, /* 0xcbfc */
            {8'h00}, /* 0xcbfb */
            {8'h00}, /* 0xcbfa */
            {8'h00}, /* 0xcbf9 */
            {8'h00}, /* 0xcbf8 */
            {8'h00}, /* 0xcbf7 */
            {8'h00}, /* 0xcbf6 */
            {8'h00}, /* 0xcbf5 */
            {8'h00}, /* 0xcbf4 */
            {8'h00}, /* 0xcbf3 */
            {8'h00}, /* 0xcbf2 */
            {8'h00}, /* 0xcbf1 */
            {8'h00}, /* 0xcbf0 */
            {8'h00}, /* 0xcbef */
            {8'h00}, /* 0xcbee */
            {8'h00}, /* 0xcbed */
            {8'h00}, /* 0xcbec */
            {8'h00}, /* 0xcbeb */
            {8'h00}, /* 0xcbea */
            {8'h00}, /* 0xcbe9 */
            {8'h00}, /* 0xcbe8 */
            {8'h00}, /* 0xcbe7 */
            {8'h00}, /* 0xcbe6 */
            {8'h00}, /* 0xcbe5 */
            {8'h00}, /* 0xcbe4 */
            {8'h00}, /* 0xcbe3 */
            {8'h00}, /* 0xcbe2 */
            {8'h00}, /* 0xcbe1 */
            {8'h00}, /* 0xcbe0 */
            {8'h00}, /* 0xcbdf */
            {8'h00}, /* 0xcbde */
            {8'h00}, /* 0xcbdd */
            {8'h00}, /* 0xcbdc */
            {8'h00}, /* 0xcbdb */
            {8'h00}, /* 0xcbda */
            {8'h00}, /* 0xcbd9 */
            {8'h00}, /* 0xcbd8 */
            {8'h00}, /* 0xcbd7 */
            {8'h00}, /* 0xcbd6 */
            {8'h00}, /* 0xcbd5 */
            {8'h00}, /* 0xcbd4 */
            {8'h00}, /* 0xcbd3 */
            {8'h00}, /* 0xcbd2 */
            {8'h00}, /* 0xcbd1 */
            {8'h00}, /* 0xcbd0 */
            {8'h00}, /* 0xcbcf */
            {8'h00}, /* 0xcbce */
            {8'h00}, /* 0xcbcd */
            {8'h00}, /* 0xcbcc */
            {8'h00}, /* 0xcbcb */
            {8'h00}, /* 0xcbca */
            {8'h00}, /* 0xcbc9 */
            {8'h00}, /* 0xcbc8 */
            {8'h00}, /* 0xcbc7 */
            {8'h00}, /* 0xcbc6 */
            {8'h00}, /* 0xcbc5 */
            {8'h00}, /* 0xcbc4 */
            {8'h00}, /* 0xcbc3 */
            {8'h00}, /* 0xcbc2 */
            {8'h00}, /* 0xcbc1 */
            {8'h00}, /* 0xcbc0 */
            {8'h00}, /* 0xcbbf */
            {8'h00}, /* 0xcbbe */
            {8'h00}, /* 0xcbbd */
            {8'h00}, /* 0xcbbc */
            {8'h00}, /* 0xcbbb */
            {8'h00}, /* 0xcbba */
            {8'h00}, /* 0xcbb9 */
            {8'h00}, /* 0xcbb8 */
            {8'h00}, /* 0xcbb7 */
            {8'h00}, /* 0xcbb6 */
            {8'h00}, /* 0xcbb5 */
            {8'h00}, /* 0xcbb4 */
            {8'h00}, /* 0xcbb3 */
            {8'h00}, /* 0xcbb2 */
            {8'h00}, /* 0xcbb1 */
            {8'h00}, /* 0xcbb0 */
            {8'h00}, /* 0xcbaf */
            {8'h00}, /* 0xcbae */
            {8'h00}, /* 0xcbad */
            {8'h00}, /* 0xcbac */
            {8'h00}, /* 0xcbab */
            {8'h00}, /* 0xcbaa */
            {8'h00}, /* 0xcba9 */
            {8'h00}, /* 0xcba8 */
            {8'h00}, /* 0xcba7 */
            {8'h00}, /* 0xcba6 */
            {8'h00}, /* 0xcba5 */
            {8'h00}, /* 0xcba4 */
            {8'h00}, /* 0xcba3 */
            {8'h00}, /* 0xcba2 */
            {8'h00}, /* 0xcba1 */
            {8'h00}, /* 0xcba0 */
            {8'h00}, /* 0xcb9f */
            {8'h00}, /* 0xcb9e */
            {8'h00}, /* 0xcb9d */
            {8'h00}, /* 0xcb9c */
            {8'h00}, /* 0xcb9b */
            {8'h00}, /* 0xcb9a */
            {8'h00}, /* 0xcb99 */
            {8'h00}, /* 0xcb98 */
            {8'h00}, /* 0xcb97 */
            {8'h00}, /* 0xcb96 */
            {8'h00}, /* 0xcb95 */
            {8'h00}, /* 0xcb94 */
            {8'h00}, /* 0xcb93 */
            {8'h00}, /* 0xcb92 */
            {8'h00}, /* 0xcb91 */
            {8'h00}, /* 0xcb90 */
            {8'h00}, /* 0xcb8f */
            {8'h00}, /* 0xcb8e */
            {8'h00}, /* 0xcb8d */
            {8'h00}, /* 0xcb8c */
            {8'h00}, /* 0xcb8b */
            {8'h00}, /* 0xcb8a */
            {8'h00}, /* 0xcb89 */
            {8'h00}, /* 0xcb88 */
            {8'h00}, /* 0xcb87 */
            {8'h00}, /* 0xcb86 */
            {8'h00}, /* 0xcb85 */
            {8'h00}, /* 0xcb84 */
            {8'h00}, /* 0xcb83 */
            {8'h00}, /* 0xcb82 */
            {8'h00}, /* 0xcb81 */
            {8'h00}, /* 0xcb80 */
            {8'h00}, /* 0xcb7f */
            {8'h00}, /* 0xcb7e */
            {8'h00}, /* 0xcb7d */
            {8'h00}, /* 0xcb7c */
            {8'h00}, /* 0xcb7b */
            {8'h00}, /* 0xcb7a */
            {8'h00}, /* 0xcb79 */
            {8'h00}, /* 0xcb78 */
            {8'h00}, /* 0xcb77 */
            {8'h00}, /* 0xcb76 */
            {8'h00}, /* 0xcb75 */
            {8'h00}, /* 0xcb74 */
            {8'h00}, /* 0xcb73 */
            {8'h00}, /* 0xcb72 */
            {8'h00}, /* 0xcb71 */
            {8'h00}, /* 0xcb70 */
            {8'h00}, /* 0xcb6f */
            {8'h00}, /* 0xcb6e */
            {8'h00}, /* 0xcb6d */
            {8'h00}, /* 0xcb6c */
            {8'h00}, /* 0xcb6b */
            {8'h00}, /* 0xcb6a */
            {8'h00}, /* 0xcb69 */
            {8'h00}, /* 0xcb68 */
            {8'h00}, /* 0xcb67 */
            {8'h00}, /* 0xcb66 */
            {8'h00}, /* 0xcb65 */
            {8'h00}, /* 0xcb64 */
            {8'h00}, /* 0xcb63 */
            {8'h00}, /* 0xcb62 */
            {8'h00}, /* 0xcb61 */
            {8'h00}, /* 0xcb60 */
            {8'h00}, /* 0xcb5f */
            {8'h00}, /* 0xcb5e */
            {8'h00}, /* 0xcb5d */
            {8'h00}, /* 0xcb5c */
            {8'h00}, /* 0xcb5b */
            {8'h00}, /* 0xcb5a */
            {8'h00}, /* 0xcb59 */
            {8'h00}, /* 0xcb58 */
            {8'h00}, /* 0xcb57 */
            {8'h00}, /* 0xcb56 */
            {8'h00}, /* 0xcb55 */
            {8'h00}, /* 0xcb54 */
            {8'h00}, /* 0xcb53 */
            {8'h00}, /* 0xcb52 */
            {8'h00}, /* 0xcb51 */
            {8'h00}, /* 0xcb50 */
            {8'h00}, /* 0xcb4f */
            {8'h00}, /* 0xcb4e */
            {8'h00}, /* 0xcb4d */
            {8'h00}, /* 0xcb4c */
            {8'h00}, /* 0xcb4b */
            {8'h00}, /* 0xcb4a */
            {8'h00}, /* 0xcb49 */
            {8'h00}, /* 0xcb48 */
            {8'h00}, /* 0xcb47 */
            {8'h00}, /* 0xcb46 */
            {8'h00}, /* 0xcb45 */
            {8'h00}, /* 0xcb44 */
            {8'h00}, /* 0xcb43 */
            {8'h00}, /* 0xcb42 */
            {8'h00}, /* 0xcb41 */
            {8'h00}, /* 0xcb40 */
            {8'h00}, /* 0xcb3f */
            {8'h00}, /* 0xcb3e */
            {8'h00}, /* 0xcb3d */
            {8'h00}, /* 0xcb3c */
            {8'h00}, /* 0xcb3b */
            {8'h00}, /* 0xcb3a */
            {8'h00}, /* 0xcb39 */
            {8'h00}, /* 0xcb38 */
            {8'h00}, /* 0xcb37 */
            {8'h00}, /* 0xcb36 */
            {8'h00}, /* 0xcb35 */
            {8'h00}, /* 0xcb34 */
            {8'h00}, /* 0xcb33 */
            {8'h00}, /* 0xcb32 */
            {8'h00}, /* 0xcb31 */
            {8'h00}, /* 0xcb30 */
            {8'h00}, /* 0xcb2f */
            {8'h00}, /* 0xcb2e */
            {8'h00}, /* 0xcb2d */
            {8'h00}, /* 0xcb2c */
            {8'h00}, /* 0xcb2b */
            {8'h00}, /* 0xcb2a */
            {8'h00}, /* 0xcb29 */
            {8'h00}, /* 0xcb28 */
            {8'h00}, /* 0xcb27 */
            {8'h00}, /* 0xcb26 */
            {8'h00}, /* 0xcb25 */
            {8'h00}, /* 0xcb24 */
            {8'h00}, /* 0xcb23 */
            {8'h00}, /* 0xcb22 */
            {8'h00}, /* 0xcb21 */
            {8'h00}, /* 0xcb20 */
            {8'h00}, /* 0xcb1f */
            {8'h00}, /* 0xcb1e */
            {8'h00}, /* 0xcb1d */
            {8'h00}, /* 0xcb1c */
            {8'h00}, /* 0xcb1b */
            {8'h00}, /* 0xcb1a */
            {8'h00}, /* 0xcb19 */
            {8'h00}, /* 0xcb18 */
            {8'h00}, /* 0xcb17 */
            {8'h00}, /* 0xcb16 */
            {8'h00}, /* 0xcb15 */
            {8'h00}, /* 0xcb14 */
            {8'h00}, /* 0xcb13 */
            {8'h00}, /* 0xcb12 */
            {8'h00}, /* 0xcb11 */
            {8'h00}, /* 0xcb10 */
            {8'h00}, /* 0xcb0f */
            {8'h00}, /* 0xcb0e */
            {8'h00}, /* 0xcb0d */
            {8'h00}, /* 0xcb0c */
            {8'h00}, /* 0xcb0b */
            {8'h00}, /* 0xcb0a */
            {8'h00}, /* 0xcb09 */
            {8'h00}, /* 0xcb08 */
            {8'h00}, /* 0xcb07 */
            {8'h00}, /* 0xcb06 */
            {8'h00}, /* 0xcb05 */
            {8'h00}, /* 0xcb04 */
            {8'h00}, /* 0xcb03 */
            {8'h00}, /* 0xcb02 */
            {8'h00}, /* 0xcb01 */
            {8'h00}, /* 0xcb00 */
            {8'h00}, /* 0xcaff */
            {8'h00}, /* 0xcafe */
            {8'h00}, /* 0xcafd */
            {8'h00}, /* 0xcafc */
            {8'h00}, /* 0xcafb */
            {8'h00}, /* 0xcafa */
            {8'h00}, /* 0xcaf9 */
            {8'h00}, /* 0xcaf8 */
            {8'h00}, /* 0xcaf7 */
            {8'h00}, /* 0xcaf6 */
            {8'h00}, /* 0xcaf5 */
            {8'h00}, /* 0xcaf4 */
            {8'h00}, /* 0xcaf3 */
            {8'h00}, /* 0xcaf2 */
            {8'h00}, /* 0xcaf1 */
            {8'h00}, /* 0xcaf0 */
            {8'h00}, /* 0xcaef */
            {8'h00}, /* 0xcaee */
            {8'h00}, /* 0xcaed */
            {8'h00}, /* 0xcaec */
            {8'h00}, /* 0xcaeb */
            {8'h00}, /* 0xcaea */
            {8'h00}, /* 0xcae9 */
            {8'h00}, /* 0xcae8 */
            {8'h00}, /* 0xcae7 */
            {8'h00}, /* 0xcae6 */
            {8'h00}, /* 0xcae5 */
            {8'h00}, /* 0xcae4 */
            {8'h00}, /* 0xcae3 */
            {8'h00}, /* 0xcae2 */
            {8'h00}, /* 0xcae1 */
            {8'h00}, /* 0xcae0 */
            {8'h00}, /* 0xcadf */
            {8'h00}, /* 0xcade */
            {8'h00}, /* 0xcadd */
            {8'h00}, /* 0xcadc */
            {8'h00}, /* 0xcadb */
            {8'h00}, /* 0xcada */
            {8'h00}, /* 0xcad9 */
            {8'h00}, /* 0xcad8 */
            {8'h00}, /* 0xcad7 */
            {8'h00}, /* 0xcad6 */
            {8'h00}, /* 0xcad5 */
            {8'h00}, /* 0xcad4 */
            {8'h00}, /* 0xcad3 */
            {8'h00}, /* 0xcad2 */
            {8'h00}, /* 0xcad1 */
            {8'h00}, /* 0xcad0 */
            {8'h00}, /* 0xcacf */
            {8'h00}, /* 0xcace */
            {8'h00}, /* 0xcacd */
            {8'h00}, /* 0xcacc */
            {8'h00}, /* 0xcacb */
            {8'h00}, /* 0xcaca */
            {8'h00}, /* 0xcac9 */
            {8'h00}, /* 0xcac8 */
            {8'h00}, /* 0xcac7 */
            {8'h00}, /* 0xcac6 */
            {8'h00}, /* 0xcac5 */
            {8'h00}, /* 0xcac4 */
            {8'h00}, /* 0xcac3 */
            {8'h00}, /* 0xcac2 */
            {8'h00}, /* 0xcac1 */
            {8'h00}, /* 0xcac0 */
            {8'h00}, /* 0xcabf */
            {8'h00}, /* 0xcabe */
            {8'h00}, /* 0xcabd */
            {8'h00}, /* 0xcabc */
            {8'h00}, /* 0xcabb */
            {8'h00}, /* 0xcaba */
            {8'h00}, /* 0xcab9 */
            {8'h00}, /* 0xcab8 */
            {8'h00}, /* 0xcab7 */
            {8'h00}, /* 0xcab6 */
            {8'h00}, /* 0xcab5 */
            {8'h00}, /* 0xcab4 */
            {8'h00}, /* 0xcab3 */
            {8'h00}, /* 0xcab2 */
            {8'h00}, /* 0xcab1 */
            {8'h00}, /* 0xcab0 */
            {8'h00}, /* 0xcaaf */
            {8'h00}, /* 0xcaae */
            {8'h00}, /* 0xcaad */
            {8'h00}, /* 0xcaac */
            {8'h00}, /* 0xcaab */
            {8'h00}, /* 0xcaaa */
            {8'h00}, /* 0xcaa9 */
            {8'h00}, /* 0xcaa8 */
            {8'h00}, /* 0xcaa7 */
            {8'h00}, /* 0xcaa6 */
            {8'h00}, /* 0xcaa5 */
            {8'h00}, /* 0xcaa4 */
            {8'h00}, /* 0xcaa3 */
            {8'h00}, /* 0xcaa2 */
            {8'h00}, /* 0xcaa1 */
            {8'h00}, /* 0xcaa0 */
            {8'h00}, /* 0xca9f */
            {8'h00}, /* 0xca9e */
            {8'h00}, /* 0xca9d */
            {8'h00}, /* 0xca9c */
            {8'h00}, /* 0xca9b */
            {8'h00}, /* 0xca9a */
            {8'h00}, /* 0xca99 */
            {8'h00}, /* 0xca98 */
            {8'h00}, /* 0xca97 */
            {8'h00}, /* 0xca96 */
            {8'h00}, /* 0xca95 */
            {8'h00}, /* 0xca94 */
            {8'h00}, /* 0xca93 */
            {8'h00}, /* 0xca92 */
            {8'h00}, /* 0xca91 */
            {8'h00}, /* 0xca90 */
            {8'h00}, /* 0xca8f */
            {8'h00}, /* 0xca8e */
            {8'h00}, /* 0xca8d */
            {8'h00}, /* 0xca8c */
            {8'h00}, /* 0xca8b */
            {8'h00}, /* 0xca8a */
            {8'h00}, /* 0xca89 */
            {8'h00}, /* 0xca88 */
            {8'h00}, /* 0xca87 */
            {8'h00}, /* 0xca86 */
            {8'h00}, /* 0xca85 */
            {8'h00}, /* 0xca84 */
            {8'h00}, /* 0xca83 */
            {8'h00}, /* 0xca82 */
            {8'h00}, /* 0xca81 */
            {8'h00}, /* 0xca80 */
            {8'h00}, /* 0xca7f */
            {8'h00}, /* 0xca7e */
            {8'h00}, /* 0xca7d */
            {8'h00}, /* 0xca7c */
            {8'h00}, /* 0xca7b */
            {8'h00}, /* 0xca7a */
            {8'h00}, /* 0xca79 */
            {8'h00}, /* 0xca78 */
            {8'h00}, /* 0xca77 */
            {8'h00}, /* 0xca76 */
            {8'h00}, /* 0xca75 */
            {8'h00}, /* 0xca74 */
            {8'h00}, /* 0xca73 */
            {8'h00}, /* 0xca72 */
            {8'h00}, /* 0xca71 */
            {8'h00}, /* 0xca70 */
            {8'h00}, /* 0xca6f */
            {8'h00}, /* 0xca6e */
            {8'h00}, /* 0xca6d */
            {8'h00}, /* 0xca6c */
            {8'h00}, /* 0xca6b */
            {8'h00}, /* 0xca6a */
            {8'h00}, /* 0xca69 */
            {8'h00}, /* 0xca68 */
            {8'h00}, /* 0xca67 */
            {8'h00}, /* 0xca66 */
            {8'h00}, /* 0xca65 */
            {8'h00}, /* 0xca64 */
            {8'h00}, /* 0xca63 */
            {8'h00}, /* 0xca62 */
            {8'h00}, /* 0xca61 */
            {8'h00}, /* 0xca60 */
            {8'h00}, /* 0xca5f */
            {8'h00}, /* 0xca5e */
            {8'h00}, /* 0xca5d */
            {8'h00}, /* 0xca5c */
            {8'h00}, /* 0xca5b */
            {8'h00}, /* 0xca5a */
            {8'h00}, /* 0xca59 */
            {8'h00}, /* 0xca58 */
            {8'h00}, /* 0xca57 */
            {8'h00}, /* 0xca56 */
            {8'h00}, /* 0xca55 */
            {8'h00}, /* 0xca54 */
            {8'h00}, /* 0xca53 */
            {8'h00}, /* 0xca52 */
            {8'h00}, /* 0xca51 */
            {8'h00}, /* 0xca50 */
            {8'h00}, /* 0xca4f */
            {8'h00}, /* 0xca4e */
            {8'h00}, /* 0xca4d */
            {8'h00}, /* 0xca4c */
            {8'h00}, /* 0xca4b */
            {8'h00}, /* 0xca4a */
            {8'h00}, /* 0xca49 */
            {8'h00}, /* 0xca48 */
            {8'h00}, /* 0xca47 */
            {8'h00}, /* 0xca46 */
            {8'h00}, /* 0xca45 */
            {8'h00}, /* 0xca44 */
            {8'h00}, /* 0xca43 */
            {8'h00}, /* 0xca42 */
            {8'h00}, /* 0xca41 */
            {8'h00}, /* 0xca40 */
            {8'h00}, /* 0xca3f */
            {8'h00}, /* 0xca3e */
            {8'h00}, /* 0xca3d */
            {8'h00}, /* 0xca3c */
            {8'h00}, /* 0xca3b */
            {8'h00}, /* 0xca3a */
            {8'h00}, /* 0xca39 */
            {8'h00}, /* 0xca38 */
            {8'h00}, /* 0xca37 */
            {8'h00}, /* 0xca36 */
            {8'h00}, /* 0xca35 */
            {8'h00}, /* 0xca34 */
            {8'h00}, /* 0xca33 */
            {8'h00}, /* 0xca32 */
            {8'h00}, /* 0xca31 */
            {8'h00}, /* 0xca30 */
            {8'h00}, /* 0xca2f */
            {8'h00}, /* 0xca2e */
            {8'h00}, /* 0xca2d */
            {8'h00}, /* 0xca2c */
            {8'h00}, /* 0xca2b */
            {8'h00}, /* 0xca2a */
            {8'h00}, /* 0xca29 */
            {8'h00}, /* 0xca28 */
            {8'h00}, /* 0xca27 */
            {8'h00}, /* 0xca26 */
            {8'h00}, /* 0xca25 */
            {8'h00}, /* 0xca24 */
            {8'h00}, /* 0xca23 */
            {8'h00}, /* 0xca22 */
            {8'h00}, /* 0xca21 */
            {8'h00}, /* 0xca20 */
            {8'h00}, /* 0xca1f */
            {8'h00}, /* 0xca1e */
            {8'h00}, /* 0xca1d */
            {8'h00}, /* 0xca1c */
            {8'h00}, /* 0xca1b */
            {8'h00}, /* 0xca1a */
            {8'h00}, /* 0xca19 */
            {8'h00}, /* 0xca18 */
            {8'h00}, /* 0xca17 */
            {8'h00}, /* 0xca16 */
            {8'h00}, /* 0xca15 */
            {8'h00}, /* 0xca14 */
            {8'h00}, /* 0xca13 */
            {8'h00}, /* 0xca12 */
            {8'h00}, /* 0xca11 */
            {8'h00}, /* 0xca10 */
            {8'h00}, /* 0xca0f */
            {8'h00}, /* 0xca0e */
            {8'h00}, /* 0xca0d */
            {8'h00}, /* 0xca0c */
            {8'h00}, /* 0xca0b */
            {8'h00}, /* 0xca0a */
            {8'h00}, /* 0xca09 */
            {8'h00}, /* 0xca08 */
            {8'h00}, /* 0xca07 */
            {8'h00}, /* 0xca06 */
            {8'h00}, /* 0xca05 */
            {8'h00}, /* 0xca04 */
            {8'h00}, /* 0xca03 */
            {8'h00}, /* 0xca02 */
            {8'h00}, /* 0xca01 */
            {8'h00}, /* 0xca00 */
            {8'h00}, /* 0xc9ff */
            {8'h00}, /* 0xc9fe */
            {8'h00}, /* 0xc9fd */
            {8'h00}, /* 0xc9fc */
            {8'h00}, /* 0xc9fb */
            {8'h00}, /* 0xc9fa */
            {8'h00}, /* 0xc9f9 */
            {8'h00}, /* 0xc9f8 */
            {8'h00}, /* 0xc9f7 */
            {8'h00}, /* 0xc9f6 */
            {8'h00}, /* 0xc9f5 */
            {8'h00}, /* 0xc9f4 */
            {8'h00}, /* 0xc9f3 */
            {8'h00}, /* 0xc9f2 */
            {8'h00}, /* 0xc9f1 */
            {8'h00}, /* 0xc9f0 */
            {8'h00}, /* 0xc9ef */
            {8'h00}, /* 0xc9ee */
            {8'h00}, /* 0xc9ed */
            {8'h00}, /* 0xc9ec */
            {8'h00}, /* 0xc9eb */
            {8'h00}, /* 0xc9ea */
            {8'h00}, /* 0xc9e9 */
            {8'h00}, /* 0xc9e8 */
            {8'h00}, /* 0xc9e7 */
            {8'h00}, /* 0xc9e6 */
            {8'h00}, /* 0xc9e5 */
            {8'h00}, /* 0xc9e4 */
            {8'h00}, /* 0xc9e3 */
            {8'h00}, /* 0xc9e2 */
            {8'h00}, /* 0xc9e1 */
            {8'h00}, /* 0xc9e0 */
            {8'h00}, /* 0xc9df */
            {8'h00}, /* 0xc9de */
            {8'h00}, /* 0xc9dd */
            {8'h00}, /* 0xc9dc */
            {8'h00}, /* 0xc9db */
            {8'h00}, /* 0xc9da */
            {8'h00}, /* 0xc9d9 */
            {8'h00}, /* 0xc9d8 */
            {8'h00}, /* 0xc9d7 */
            {8'h00}, /* 0xc9d6 */
            {8'h00}, /* 0xc9d5 */
            {8'h00}, /* 0xc9d4 */
            {8'h00}, /* 0xc9d3 */
            {8'h00}, /* 0xc9d2 */
            {8'h00}, /* 0xc9d1 */
            {8'h00}, /* 0xc9d0 */
            {8'h00}, /* 0xc9cf */
            {8'h00}, /* 0xc9ce */
            {8'h00}, /* 0xc9cd */
            {8'h00}, /* 0xc9cc */
            {8'h00}, /* 0xc9cb */
            {8'h00}, /* 0xc9ca */
            {8'h00}, /* 0xc9c9 */
            {8'h00}, /* 0xc9c8 */
            {8'h00}, /* 0xc9c7 */
            {8'h00}, /* 0xc9c6 */
            {8'h00}, /* 0xc9c5 */
            {8'h00}, /* 0xc9c4 */
            {8'h00}, /* 0xc9c3 */
            {8'h00}, /* 0xc9c2 */
            {8'h00}, /* 0xc9c1 */
            {8'h00}, /* 0xc9c0 */
            {8'h00}, /* 0xc9bf */
            {8'h00}, /* 0xc9be */
            {8'h00}, /* 0xc9bd */
            {8'h00}, /* 0xc9bc */
            {8'h00}, /* 0xc9bb */
            {8'h00}, /* 0xc9ba */
            {8'h00}, /* 0xc9b9 */
            {8'h00}, /* 0xc9b8 */
            {8'h00}, /* 0xc9b7 */
            {8'h00}, /* 0xc9b6 */
            {8'h00}, /* 0xc9b5 */
            {8'h00}, /* 0xc9b4 */
            {8'h00}, /* 0xc9b3 */
            {8'h00}, /* 0xc9b2 */
            {8'h00}, /* 0xc9b1 */
            {8'h00}, /* 0xc9b0 */
            {8'h00}, /* 0xc9af */
            {8'h00}, /* 0xc9ae */
            {8'h00}, /* 0xc9ad */
            {8'h00}, /* 0xc9ac */
            {8'h00}, /* 0xc9ab */
            {8'h00}, /* 0xc9aa */
            {8'h00}, /* 0xc9a9 */
            {8'h00}, /* 0xc9a8 */
            {8'h00}, /* 0xc9a7 */
            {8'h00}, /* 0xc9a6 */
            {8'h00}, /* 0xc9a5 */
            {8'h00}, /* 0xc9a4 */
            {8'h00}, /* 0xc9a3 */
            {8'h00}, /* 0xc9a2 */
            {8'h00}, /* 0xc9a1 */
            {8'h00}, /* 0xc9a0 */
            {8'h00}, /* 0xc99f */
            {8'h00}, /* 0xc99e */
            {8'h00}, /* 0xc99d */
            {8'h00}, /* 0xc99c */
            {8'h00}, /* 0xc99b */
            {8'h00}, /* 0xc99a */
            {8'h00}, /* 0xc999 */
            {8'h00}, /* 0xc998 */
            {8'h00}, /* 0xc997 */
            {8'h00}, /* 0xc996 */
            {8'h00}, /* 0xc995 */
            {8'h00}, /* 0xc994 */
            {8'h00}, /* 0xc993 */
            {8'h00}, /* 0xc992 */
            {8'h00}, /* 0xc991 */
            {8'h00}, /* 0xc990 */
            {8'h00}, /* 0xc98f */
            {8'h00}, /* 0xc98e */
            {8'h00}, /* 0xc98d */
            {8'h00}, /* 0xc98c */
            {8'h00}, /* 0xc98b */
            {8'h00}, /* 0xc98a */
            {8'h00}, /* 0xc989 */
            {8'h00}, /* 0xc988 */
            {8'h00}, /* 0xc987 */
            {8'h00}, /* 0xc986 */
            {8'h00}, /* 0xc985 */
            {8'h00}, /* 0xc984 */
            {8'h00}, /* 0xc983 */
            {8'h00}, /* 0xc982 */
            {8'h00}, /* 0xc981 */
            {8'h00}, /* 0xc980 */
            {8'h00}, /* 0xc97f */
            {8'h00}, /* 0xc97e */
            {8'h00}, /* 0xc97d */
            {8'h00}, /* 0xc97c */
            {8'h00}, /* 0xc97b */
            {8'h00}, /* 0xc97a */
            {8'h00}, /* 0xc979 */
            {8'h00}, /* 0xc978 */
            {8'h00}, /* 0xc977 */
            {8'h00}, /* 0xc976 */
            {8'h00}, /* 0xc975 */
            {8'h00}, /* 0xc974 */
            {8'h00}, /* 0xc973 */
            {8'h00}, /* 0xc972 */
            {8'h00}, /* 0xc971 */
            {8'h00}, /* 0xc970 */
            {8'h00}, /* 0xc96f */
            {8'h00}, /* 0xc96e */
            {8'h00}, /* 0xc96d */
            {8'h00}, /* 0xc96c */
            {8'h00}, /* 0xc96b */
            {8'h00}, /* 0xc96a */
            {8'h00}, /* 0xc969 */
            {8'h00}, /* 0xc968 */
            {8'h00}, /* 0xc967 */
            {8'h00}, /* 0xc966 */
            {8'h00}, /* 0xc965 */
            {8'h00}, /* 0xc964 */
            {8'h00}, /* 0xc963 */
            {8'h00}, /* 0xc962 */
            {8'h00}, /* 0xc961 */
            {8'h00}, /* 0xc960 */
            {8'h00}, /* 0xc95f */
            {8'h00}, /* 0xc95e */
            {8'h00}, /* 0xc95d */
            {8'h00}, /* 0xc95c */
            {8'h00}, /* 0xc95b */
            {8'h00}, /* 0xc95a */
            {8'h00}, /* 0xc959 */
            {8'h00}, /* 0xc958 */
            {8'h00}, /* 0xc957 */
            {8'h00}, /* 0xc956 */
            {8'h00}, /* 0xc955 */
            {8'h00}, /* 0xc954 */
            {8'h00}, /* 0xc953 */
            {8'h00}, /* 0xc952 */
            {8'h00}, /* 0xc951 */
            {8'h00}, /* 0xc950 */
            {8'h00}, /* 0xc94f */
            {8'h00}, /* 0xc94e */
            {8'h00}, /* 0xc94d */
            {8'h00}, /* 0xc94c */
            {8'h00}, /* 0xc94b */
            {8'h00}, /* 0xc94a */
            {8'h00}, /* 0xc949 */
            {8'h00}, /* 0xc948 */
            {8'h00}, /* 0xc947 */
            {8'h00}, /* 0xc946 */
            {8'h00}, /* 0xc945 */
            {8'h00}, /* 0xc944 */
            {8'h00}, /* 0xc943 */
            {8'h00}, /* 0xc942 */
            {8'h00}, /* 0xc941 */
            {8'h00}, /* 0xc940 */
            {8'h00}, /* 0xc93f */
            {8'h00}, /* 0xc93e */
            {8'h00}, /* 0xc93d */
            {8'h00}, /* 0xc93c */
            {8'h00}, /* 0xc93b */
            {8'h00}, /* 0xc93a */
            {8'h00}, /* 0xc939 */
            {8'h00}, /* 0xc938 */
            {8'h00}, /* 0xc937 */
            {8'h00}, /* 0xc936 */
            {8'h00}, /* 0xc935 */
            {8'h00}, /* 0xc934 */
            {8'h00}, /* 0xc933 */
            {8'h00}, /* 0xc932 */
            {8'h00}, /* 0xc931 */
            {8'h00}, /* 0xc930 */
            {8'h00}, /* 0xc92f */
            {8'h00}, /* 0xc92e */
            {8'h00}, /* 0xc92d */
            {8'h00}, /* 0xc92c */
            {8'h00}, /* 0xc92b */
            {8'h00}, /* 0xc92a */
            {8'h00}, /* 0xc929 */
            {8'h00}, /* 0xc928 */
            {8'h00}, /* 0xc927 */
            {8'h00}, /* 0xc926 */
            {8'h00}, /* 0xc925 */
            {8'h00}, /* 0xc924 */
            {8'h00}, /* 0xc923 */
            {8'h00}, /* 0xc922 */
            {8'h00}, /* 0xc921 */
            {8'h00}, /* 0xc920 */
            {8'h00}, /* 0xc91f */
            {8'h00}, /* 0xc91e */
            {8'h00}, /* 0xc91d */
            {8'h00}, /* 0xc91c */
            {8'h00}, /* 0xc91b */
            {8'h00}, /* 0xc91a */
            {8'h00}, /* 0xc919 */
            {8'h00}, /* 0xc918 */
            {8'h00}, /* 0xc917 */
            {8'h00}, /* 0xc916 */
            {8'h00}, /* 0xc915 */
            {8'h00}, /* 0xc914 */
            {8'h00}, /* 0xc913 */
            {8'h00}, /* 0xc912 */
            {8'h00}, /* 0xc911 */
            {8'h00}, /* 0xc910 */
            {8'h00}, /* 0xc90f */
            {8'h00}, /* 0xc90e */
            {8'h00}, /* 0xc90d */
            {8'h00}, /* 0xc90c */
            {8'h00}, /* 0xc90b */
            {8'h00}, /* 0xc90a */
            {8'h00}, /* 0xc909 */
            {8'h00}, /* 0xc908 */
            {8'h00}, /* 0xc907 */
            {8'h00}, /* 0xc906 */
            {8'h00}, /* 0xc905 */
            {8'h00}, /* 0xc904 */
            {8'h00}, /* 0xc903 */
            {8'h00}, /* 0xc902 */
            {8'h00}, /* 0xc901 */
            {8'h00}, /* 0xc900 */
            {8'h00}, /* 0xc8ff */
            {8'h00}, /* 0xc8fe */
            {8'h00}, /* 0xc8fd */
            {8'h00}, /* 0xc8fc */
            {8'h00}, /* 0xc8fb */
            {8'h00}, /* 0xc8fa */
            {8'h00}, /* 0xc8f9 */
            {8'h00}, /* 0xc8f8 */
            {8'h00}, /* 0xc8f7 */
            {8'h00}, /* 0xc8f6 */
            {8'h00}, /* 0xc8f5 */
            {8'h00}, /* 0xc8f4 */
            {8'h00}, /* 0xc8f3 */
            {8'h00}, /* 0xc8f2 */
            {8'h00}, /* 0xc8f1 */
            {8'h00}, /* 0xc8f0 */
            {8'h00}, /* 0xc8ef */
            {8'h00}, /* 0xc8ee */
            {8'h00}, /* 0xc8ed */
            {8'h00}, /* 0xc8ec */
            {8'h00}, /* 0xc8eb */
            {8'h00}, /* 0xc8ea */
            {8'h00}, /* 0xc8e9 */
            {8'h00}, /* 0xc8e8 */
            {8'h00}, /* 0xc8e7 */
            {8'h00}, /* 0xc8e6 */
            {8'h00}, /* 0xc8e5 */
            {8'h00}, /* 0xc8e4 */
            {8'h00}, /* 0xc8e3 */
            {8'h00}, /* 0xc8e2 */
            {8'h00}, /* 0xc8e1 */
            {8'h00}, /* 0xc8e0 */
            {8'h00}, /* 0xc8df */
            {8'h00}, /* 0xc8de */
            {8'h00}, /* 0xc8dd */
            {8'h00}, /* 0xc8dc */
            {8'h00}, /* 0xc8db */
            {8'h00}, /* 0xc8da */
            {8'h00}, /* 0xc8d9 */
            {8'h00}, /* 0xc8d8 */
            {8'h00}, /* 0xc8d7 */
            {8'h00}, /* 0xc8d6 */
            {8'h00}, /* 0xc8d5 */
            {8'h00}, /* 0xc8d4 */
            {8'h00}, /* 0xc8d3 */
            {8'h00}, /* 0xc8d2 */
            {8'h00}, /* 0xc8d1 */
            {8'h00}, /* 0xc8d0 */
            {8'h00}, /* 0xc8cf */
            {8'h00}, /* 0xc8ce */
            {8'h00}, /* 0xc8cd */
            {8'h00}, /* 0xc8cc */
            {8'h00}, /* 0xc8cb */
            {8'h00}, /* 0xc8ca */
            {8'h00}, /* 0xc8c9 */
            {8'h00}, /* 0xc8c8 */
            {8'h00}, /* 0xc8c7 */
            {8'h00}, /* 0xc8c6 */
            {8'h00}, /* 0xc8c5 */
            {8'h00}, /* 0xc8c4 */
            {8'h00}, /* 0xc8c3 */
            {8'h00}, /* 0xc8c2 */
            {8'h00}, /* 0xc8c1 */
            {8'h00}, /* 0xc8c0 */
            {8'h00}, /* 0xc8bf */
            {8'h00}, /* 0xc8be */
            {8'h00}, /* 0xc8bd */
            {8'h00}, /* 0xc8bc */
            {8'h00}, /* 0xc8bb */
            {8'h00}, /* 0xc8ba */
            {8'h00}, /* 0xc8b9 */
            {8'h00}, /* 0xc8b8 */
            {8'h00}, /* 0xc8b7 */
            {8'h00}, /* 0xc8b6 */
            {8'h00}, /* 0xc8b5 */
            {8'h00}, /* 0xc8b4 */
            {8'h00}, /* 0xc8b3 */
            {8'h00}, /* 0xc8b2 */
            {8'h00}, /* 0xc8b1 */
            {8'h00}, /* 0xc8b0 */
            {8'h00}, /* 0xc8af */
            {8'h00}, /* 0xc8ae */
            {8'h00}, /* 0xc8ad */
            {8'h00}, /* 0xc8ac */
            {8'h00}, /* 0xc8ab */
            {8'h00}, /* 0xc8aa */
            {8'h00}, /* 0xc8a9 */
            {8'h00}, /* 0xc8a8 */
            {8'h00}, /* 0xc8a7 */
            {8'h00}, /* 0xc8a6 */
            {8'h00}, /* 0xc8a5 */
            {8'h00}, /* 0xc8a4 */
            {8'h00}, /* 0xc8a3 */
            {8'h00}, /* 0xc8a2 */
            {8'h00}, /* 0xc8a1 */
            {8'h00}, /* 0xc8a0 */
            {8'h00}, /* 0xc89f */
            {8'h00}, /* 0xc89e */
            {8'h00}, /* 0xc89d */
            {8'h00}, /* 0xc89c */
            {8'h00}, /* 0xc89b */
            {8'h00}, /* 0xc89a */
            {8'h00}, /* 0xc899 */
            {8'h00}, /* 0xc898 */
            {8'h00}, /* 0xc897 */
            {8'h00}, /* 0xc896 */
            {8'h00}, /* 0xc895 */
            {8'h00}, /* 0xc894 */
            {8'h00}, /* 0xc893 */
            {8'h00}, /* 0xc892 */
            {8'h00}, /* 0xc891 */
            {8'h00}, /* 0xc890 */
            {8'h00}, /* 0xc88f */
            {8'h00}, /* 0xc88e */
            {8'h00}, /* 0xc88d */
            {8'h00}, /* 0xc88c */
            {8'h00}, /* 0xc88b */
            {8'h00}, /* 0xc88a */
            {8'h00}, /* 0xc889 */
            {8'h00}, /* 0xc888 */
            {8'h00}, /* 0xc887 */
            {8'h00}, /* 0xc886 */
            {8'h00}, /* 0xc885 */
            {8'h00}, /* 0xc884 */
            {8'h00}, /* 0xc883 */
            {8'h00}, /* 0xc882 */
            {8'h00}, /* 0xc881 */
            {8'h00}, /* 0xc880 */
            {8'h00}, /* 0xc87f */
            {8'h00}, /* 0xc87e */
            {8'h00}, /* 0xc87d */
            {8'h00}, /* 0xc87c */
            {8'h00}, /* 0xc87b */
            {8'h00}, /* 0xc87a */
            {8'h00}, /* 0xc879 */
            {8'h00}, /* 0xc878 */
            {8'h00}, /* 0xc877 */
            {8'h00}, /* 0xc876 */
            {8'h00}, /* 0xc875 */
            {8'h00}, /* 0xc874 */
            {8'h00}, /* 0xc873 */
            {8'h00}, /* 0xc872 */
            {8'h00}, /* 0xc871 */
            {8'h00}, /* 0xc870 */
            {8'h00}, /* 0xc86f */
            {8'h00}, /* 0xc86e */
            {8'h00}, /* 0xc86d */
            {8'h00}, /* 0xc86c */
            {8'h00}, /* 0xc86b */
            {8'h00}, /* 0xc86a */
            {8'h00}, /* 0xc869 */
            {8'h00}, /* 0xc868 */
            {8'h00}, /* 0xc867 */
            {8'h00}, /* 0xc866 */
            {8'h00}, /* 0xc865 */
            {8'h00}, /* 0xc864 */
            {8'h00}, /* 0xc863 */
            {8'h00}, /* 0xc862 */
            {8'h00}, /* 0xc861 */
            {8'h00}, /* 0xc860 */
            {8'h00}, /* 0xc85f */
            {8'h00}, /* 0xc85e */
            {8'h00}, /* 0xc85d */
            {8'h00}, /* 0xc85c */
            {8'h00}, /* 0xc85b */
            {8'h00}, /* 0xc85a */
            {8'h00}, /* 0xc859 */
            {8'h00}, /* 0xc858 */
            {8'h00}, /* 0xc857 */
            {8'h00}, /* 0xc856 */
            {8'h00}, /* 0xc855 */
            {8'h00}, /* 0xc854 */
            {8'h00}, /* 0xc853 */
            {8'h00}, /* 0xc852 */
            {8'h00}, /* 0xc851 */
            {8'h00}, /* 0xc850 */
            {8'h00}, /* 0xc84f */
            {8'h00}, /* 0xc84e */
            {8'h00}, /* 0xc84d */
            {8'h00}, /* 0xc84c */
            {8'h00}, /* 0xc84b */
            {8'h00}, /* 0xc84a */
            {8'h00}, /* 0xc849 */
            {8'h00}, /* 0xc848 */
            {8'h00}, /* 0xc847 */
            {8'h00}, /* 0xc846 */
            {8'h00}, /* 0xc845 */
            {8'h00}, /* 0xc844 */
            {8'h00}, /* 0xc843 */
            {8'h00}, /* 0xc842 */
            {8'h00}, /* 0xc841 */
            {8'h00}, /* 0xc840 */
            {8'h00}, /* 0xc83f */
            {8'h00}, /* 0xc83e */
            {8'h00}, /* 0xc83d */
            {8'h00}, /* 0xc83c */
            {8'h00}, /* 0xc83b */
            {8'h00}, /* 0xc83a */
            {8'h00}, /* 0xc839 */
            {8'h00}, /* 0xc838 */
            {8'h00}, /* 0xc837 */
            {8'h00}, /* 0xc836 */
            {8'h00}, /* 0xc835 */
            {8'h00}, /* 0xc834 */
            {8'h00}, /* 0xc833 */
            {8'h00}, /* 0xc832 */
            {8'h00}, /* 0xc831 */
            {8'h00}, /* 0xc830 */
            {8'h00}, /* 0xc82f */
            {8'h00}, /* 0xc82e */
            {8'h00}, /* 0xc82d */
            {8'h00}, /* 0xc82c */
            {8'h00}, /* 0xc82b */
            {8'h00}, /* 0xc82a */
            {8'h00}, /* 0xc829 */
            {8'h00}, /* 0xc828 */
            {8'h00}, /* 0xc827 */
            {8'h00}, /* 0xc826 */
            {8'h00}, /* 0xc825 */
            {8'h00}, /* 0xc824 */
            {8'h00}, /* 0xc823 */
            {8'h00}, /* 0xc822 */
            {8'h00}, /* 0xc821 */
            {8'h00}, /* 0xc820 */
            {8'h00}, /* 0xc81f */
            {8'h00}, /* 0xc81e */
            {8'h00}, /* 0xc81d */
            {8'h00}, /* 0xc81c */
            {8'h00}, /* 0xc81b */
            {8'h00}, /* 0xc81a */
            {8'h00}, /* 0xc819 */
            {8'h00}, /* 0xc818 */
            {8'h00}, /* 0xc817 */
            {8'h00}, /* 0xc816 */
            {8'h00}, /* 0xc815 */
            {8'h00}, /* 0xc814 */
            {8'h00}, /* 0xc813 */
            {8'h00}, /* 0xc812 */
            {8'h00}, /* 0xc811 */
            {8'h00}, /* 0xc810 */
            {8'h00}, /* 0xc80f */
            {8'h00}, /* 0xc80e */
            {8'h00}, /* 0xc80d */
            {8'h00}, /* 0xc80c */
            {8'h00}, /* 0xc80b */
            {8'h00}, /* 0xc80a */
            {8'h00}, /* 0xc809 */
            {8'h00}, /* 0xc808 */
            {8'h00}, /* 0xc807 */
            {8'h00}, /* 0xc806 */
            {8'h00}, /* 0xc805 */
            {8'h00}, /* 0xc804 */
            {8'h00}, /* 0xc803 */
            {8'h00}, /* 0xc802 */
            {8'h00}, /* 0xc801 */
            {8'h00}, /* 0xc800 */
            {8'h00}, /* 0xc7ff */
            {8'h00}, /* 0xc7fe */
            {8'h00}, /* 0xc7fd */
            {8'h00}, /* 0xc7fc */
            {8'h00}, /* 0xc7fb */
            {8'h00}, /* 0xc7fa */
            {8'h00}, /* 0xc7f9 */
            {8'h00}, /* 0xc7f8 */
            {8'h00}, /* 0xc7f7 */
            {8'h00}, /* 0xc7f6 */
            {8'h00}, /* 0xc7f5 */
            {8'h00}, /* 0xc7f4 */
            {8'h00}, /* 0xc7f3 */
            {8'h00}, /* 0xc7f2 */
            {8'h00}, /* 0xc7f1 */
            {8'h00}, /* 0xc7f0 */
            {8'h00}, /* 0xc7ef */
            {8'h00}, /* 0xc7ee */
            {8'h00}, /* 0xc7ed */
            {8'h00}, /* 0xc7ec */
            {8'h00}, /* 0xc7eb */
            {8'h00}, /* 0xc7ea */
            {8'h00}, /* 0xc7e9 */
            {8'h00}, /* 0xc7e8 */
            {8'h00}, /* 0xc7e7 */
            {8'h00}, /* 0xc7e6 */
            {8'h00}, /* 0xc7e5 */
            {8'h00}, /* 0xc7e4 */
            {8'h00}, /* 0xc7e3 */
            {8'h00}, /* 0xc7e2 */
            {8'h00}, /* 0xc7e1 */
            {8'h00}, /* 0xc7e0 */
            {8'h00}, /* 0xc7df */
            {8'h00}, /* 0xc7de */
            {8'h00}, /* 0xc7dd */
            {8'h00}, /* 0xc7dc */
            {8'h00}, /* 0xc7db */
            {8'h00}, /* 0xc7da */
            {8'h00}, /* 0xc7d9 */
            {8'h00}, /* 0xc7d8 */
            {8'h00}, /* 0xc7d7 */
            {8'h00}, /* 0xc7d6 */
            {8'h00}, /* 0xc7d5 */
            {8'h00}, /* 0xc7d4 */
            {8'h00}, /* 0xc7d3 */
            {8'h00}, /* 0xc7d2 */
            {8'h00}, /* 0xc7d1 */
            {8'h00}, /* 0xc7d0 */
            {8'h00}, /* 0xc7cf */
            {8'h00}, /* 0xc7ce */
            {8'h00}, /* 0xc7cd */
            {8'h00}, /* 0xc7cc */
            {8'h00}, /* 0xc7cb */
            {8'h00}, /* 0xc7ca */
            {8'h00}, /* 0xc7c9 */
            {8'h00}, /* 0xc7c8 */
            {8'h00}, /* 0xc7c7 */
            {8'h00}, /* 0xc7c6 */
            {8'h00}, /* 0xc7c5 */
            {8'h00}, /* 0xc7c4 */
            {8'h00}, /* 0xc7c3 */
            {8'h00}, /* 0xc7c2 */
            {8'h00}, /* 0xc7c1 */
            {8'h00}, /* 0xc7c0 */
            {8'h00}, /* 0xc7bf */
            {8'h00}, /* 0xc7be */
            {8'h00}, /* 0xc7bd */
            {8'h00}, /* 0xc7bc */
            {8'h00}, /* 0xc7bb */
            {8'h00}, /* 0xc7ba */
            {8'h00}, /* 0xc7b9 */
            {8'h00}, /* 0xc7b8 */
            {8'h00}, /* 0xc7b7 */
            {8'h00}, /* 0xc7b6 */
            {8'h00}, /* 0xc7b5 */
            {8'h00}, /* 0xc7b4 */
            {8'h00}, /* 0xc7b3 */
            {8'h00}, /* 0xc7b2 */
            {8'h00}, /* 0xc7b1 */
            {8'h00}, /* 0xc7b0 */
            {8'h00}, /* 0xc7af */
            {8'h00}, /* 0xc7ae */
            {8'h00}, /* 0xc7ad */
            {8'h00}, /* 0xc7ac */
            {8'h00}, /* 0xc7ab */
            {8'h00}, /* 0xc7aa */
            {8'h00}, /* 0xc7a9 */
            {8'h00}, /* 0xc7a8 */
            {8'h00}, /* 0xc7a7 */
            {8'h00}, /* 0xc7a6 */
            {8'h00}, /* 0xc7a5 */
            {8'h00}, /* 0xc7a4 */
            {8'h00}, /* 0xc7a3 */
            {8'h00}, /* 0xc7a2 */
            {8'h00}, /* 0xc7a1 */
            {8'h00}, /* 0xc7a0 */
            {8'h00}, /* 0xc79f */
            {8'h00}, /* 0xc79e */
            {8'h00}, /* 0xc79d */
            {8'h00}, /* 0xc79c */
            {8'h00}, /* 0xc79b */
            {8'h00}, /* 0xc79a */
            {8'h00}, /* 0xc799 */
            {8'h00}, /* 0xc798 */
            {8'h00}, /* 0xc797 */
            {8'h00}, /* 0xc796 */
            {8'h00}, /* 0xc795 */
            {8'h00}, /* 0xc794 */
            {8'h00}, /* 0xc793 */
            {8'h00}, /* 0xc792 */
            {8'h00}, /* 0xc791 */
            {8'h00}, /* 0xc790 */
            {8'h00}, /* 0xc78f */
            {8'h00}, /* 0xc78e */
            {8'h00}, /* 0xc78d */
            {8'h00}, /* 0xc78c */
            {8'h00}, /* 0xc78b */
            {8'h00}, /* 0xc78a */
            {8'h00}, /* 0xc789 */
            {8'h00}, /* 0xc788 */
            {8'h00}, /* 0xc787 */
            {8'h00}, /* 0xc786 */
            {8'h00}, /* 0xc785 */
            {8'h00}, /* 0xc784 */
            {8'h00}, /* 0xc783 */
            {8'h00}, /* 0xc782 */
            {8'h00}, /* 0xc781 */
            {8'h00}, /* 0xc780 */
            {8'h00}, /* 0xc77f */
            {8'h00}, /* 0xc77e */
            {8'h00}, /* 0xc77d */
            {8'h00}, /* 0xc77c */
            {8'h00}, /* 0xc77b */
            {8'h00}, /* 0xc77a */
            {8'h00}, /* 0xc779 */
            {8'h00}, /* 0xc778 */
            {8'h00}, /* 0xc777 */
            {8'h00}, /* 0xc776 */
            {8'h00}, /* 0xc775 */
            {8'h00}, /* 0xc774 */
            {8'h00}, /* 0xc773 */
            {8'h00}, /* 0xc772 */
            {8'h00}, /* 0xc771 */
            {8'h00}, /* 0xc770 */
            {8'h00}, /* 0xc76f */
            {8'h00}, /* 0xc76e */
            {8'h00}, /* 0xc76d */
            {8'h00}, /* 0xc76c */
            {8'h00}, /* 0xc76b */
            {8'h00}, /* 0xc76a */
            {8'h00}, /* 0xc769 */
            {8'h00}, /* 0xc768 */
            {8'h00}, /* 0xc767 */
            {8'h00}, /* 0xc766 */
            {8'h00}, /* 0xc765 */
            {8'h00}, /* 0xc764 */
            {8'h00}, /* 0xc763 */
            {8'h00}, /* 0xc762 */
            {8'h00}, /* 0xc761 */
            {8'h00}, /* 0xc760 */
            {8'h00}, /* 0xc75f */
            {8'h00}, /* 0xc75e */
            {8'h00}, /* 0xc75d */
            {8'h00}, /* 0xc75c */
            {8'h00}, /* 0xc75b */
            {8'h00}, /* 0xc75a */
            {8'h00}, /* 0xc759 */
            {8'h00}, /* 0xc758 */
            {8'h00}, /* 0xc757 */
            {8'h00}, /* 0xc756 */
            {8'h00}, /* 0xc755 */
            {8'h00}, /* 0xc754 */
            {8'h00}, /* 0xc753 */
            {8'h00}, /* 0xc752 */
            {8'h00}, /* 0xc751 */
            {8'h00}, /* 0xc750 */
            {8'h00}, /* 0xc74f */
            {8'h00}, /* 0xc74e */
            {8'h00}, /* 0xc74d */
            {8'h00}, /* 0xc74c */
            {8'h00}, /* 0xc74b */
            {8'h00}, /* 0xc74a */
            {8'h00}, /* 0xc749 */
            {8'h00}, /* 0xc748 */
            {8'h00}, /* 0xc747 */
            {8'h00}, /* 0xc746 */
            {8'h00}, /* 0xc745 */
            {8'h00}, /* 0xc744 */
            {8'h00}, /* 0xc743 */
            {8'h00}, /* 0xc742 */
            {8'h00}, /* 0xc741 */
            {8'h00}, /* 0xc740 */
            {8'h00}, /* 0xc73f */
            {8'h00}, /* 0xc73e */
            {8'h00}, /* 0xc73d */
            {8'h00}, /* 0xc73c */
            {8'h00}, /* 0xc73b */
            {8'h00}, /* 0xc73a */
            {8'h00}, /* 0xc739 */
            {8'h00}, /* 0xc738 */
            {8'h00}, /* 0xc737 */
            {8'h00}, /* 0xc736 */
            {8'h00}, /* 0xc735 */
            {8'h00}, /* 0xc734 */
            {8'h00}, /* 0xc733 */
            {8'h00}, /* 0xc732 */
            {8'h00}, /* 0xc731 */
            {8'h00}, /* 0xc730 */
            {8'h00}, /* 0xc72f */
            {8'h00}, /* 0xc72e */
            {8'h00}, /* 0xc72d */
            {8'h00}, /* 0xc72c */
            {8'h00}, /* 0xc72b */
            {8'h00}, /* 0xc72a */
            {8'h00}, /* 0xc729 */
            {8'h00}, /* 0xc728 */
            {8'h00}, /* 0xc727 */
            {8'h00}, /* 0xc726 */
            {8'h00}, /* 0xc725 */
            {8'h00}, /* 0xc724 */
            {8'h00}, /* 0xc723 */
            {8'h00}, /* 0xc722 */
            {8'h00}, /* 0xc721 */
            {8'h00}, /* 0xc720 */
            {8'h00}, /* 0xc71f */
            {8'h00}, /* 0xc71e */
            {8'h00}, /* 0xc71d */
            {8'h00}, /* 0xc71c */
            {8'h00}, /* 0xc71b */
            {8'h00}, /* 0xc71a */
            {8'h00}, /* 0xc719 */
            {8'h00}, /* 0xc718 */
            {8'h00}, /* 0xc717 */
            {8'h00}, /* 0xc716 */
            {8'h00}, /* 0xc715 */
            {8'h00}, /* 0xc714 */
            {8'h00}, /* 0xc713 */
            {8'h00}, /* 0xc712 */
            {8'h00}, /* 0xc711 */
            {8'h00}, /* 0xc710 */
            {8'h00}, /* 0xc70f */
            {8'h00}, /* 0xc70e */
            {8'h00}, /* 0xc70d */
            {8'h00}, /* 0xc70c */
            {8'h00}, /* 0xc70b */
            {8'h00}, /* 0xc70a */
            {8'h00}, /* 0xc709 */
            {8'h00}, /* 0xc708 */
            {8'h00}, /* 0xc707 */
            {8'h00}, /* 0xc706 */
            {8'h00}, /* 0xc705 */
            {8'h00}, /* 0xc704 */
            {8'h00}, /* 0xc703 */
            {8'h00}, /* 0xc702 */
            {8'h00}, /* 0xc701 */
            {8'h00}, /* 0xc700 */
            {8'h00}, /* 0xc6ff */
            {8'h00}, /* 0xc6fe */
            {8'h00}, /* 0xc6fd */
            {8'h00}, /* 0xc6fc */
            {8'h00}, /* 0xc6fb */
            {8'h00}, /* 0xc6fa */
            {8'h00}, /* 0xc6f9 */
            {8'h00}, /* 0xc6f8 */
            {8'h00}, /* 0xc6f7 */
            {8'h00}, /* 0xc6f6 */
            {8'h00}, /* 0xc6f5 */
            {8'h00}, /* 0xc6f4 */
            {8'h00}, /* 0xc6f3 */
            {8'h00}, /* 0xc6f2 */
            {8'h00}, /* 0xc6f1 */
            {8'h00}, /* 0xc6f0 */
            {8'h00}, /* 0xc6ef */
            {8'h00}, /* 0xc6ee */
            {8'h00}, /* 0xc6ed */
            {8'h00}, /* 0xc6ec */
            {8'h00}, /* 0xc6eb */
            {8'h00}, /* 0xc6ea */
            {8'h00}, /* 0xc6e9 */
            {8'h00}, /* 0xc6e8 */
            {8'h00}, /* 0xc6e7 */
            {8'h00}, /* 0xc6e6 */
            {8'h00}, /* 0xc6e5 */
            {8'h00}, /* 0xc6e4 */
            {8'h00}, /* 0xc6e3 */
            {8'h00}, /* 0xc6e2 */
            {8'h00}, /* 0xc6e1 */
            {8'h00}, /* 0xc6e0 */
            {8'h00}, /* 0xc6df */
            {8'h00}, /* 0xc6de */
            {8'h00}, /* 0xc6dd */
            {8'h00}, /* 0xc6dc */
            {8'h00}, /* 0xc6db */
            {8'h00}, /* 0xc6da */
            {8'h00}, /* 0xc6d9 */
            {8'h00}, /* 0xc6d8 */
            {8'h00}, /* 0xc6d7 */
            {8'h00}, /* 0xc6d6 */
            {8'h00}, /* 0xc6d5 */
            {8'h00}, /* 0xc6d4 */
            {8'h00}, /* 0xc6d3 */
            {8'h00}, /* 0xc6d2 */
            {8'h00}, /* 0xc6d1 */
            {8'h00}, /* 0xc6d0 */
            {8'h00}, /* 0xc6cf */
            {8'h00}, /* 0xc6ce */
            {8'h00}, /* 0xc6cd */
            {8'h00}, /* 0xc6cc */
            {8'h00}, /* 0xc6cb */
            {8'h00}, /* 0xc6ca */
            {8'h00}, /* 0xc6c9 */
            {8'h00}, /* 0xc6c8 */
            {8'h00}, /* 0xc6c7 */
            {8'h00}, /* 0xc6c6 */
            {8'h00}, /* 0xc6c5 */
            {8'h00}, /* 0xc6c4 */
            {8'h00}, /* 0xc6c3 */
            {8'h00}, /* 0xc6c2 */
            {8'h00}, /* 0xc6c1 */
            {8'h00}, /* 0xc6c0 */
            {8'h00}, /* 0xc6bf */
            {8'h00}, /* 0xc6be */
            {8'h00}, /* 0xc6bd */
            {8'h00}, /* 0xc6bc */
            {8'h00}, /* 0xc6bb */
            {8'h00}, /* 0xc6ba */
            {8'h00}, /* 0xc6b9 */
            {8'h00}, /* 0xc6b8 */
            {8'h00}, /* 0xc6b7 */
            {8'h00}, /* 0xc6b6 */
            {8'h00}, /* 0xc6b5 */
            {8'h00}, /* 0xc6b4 */
            {8'h00}, /* 0xc6b3 */
            {8'h00}, /* 0xc6b2 */
            {8'h00}, /* 0xc6b1 */
            {8'h00}, /* 0xc6b0 */
            {8'h00}, /* 0xc6af */
            {8'h00}, /* 0xc6ae */
            {8'h00}, /* 0xc6ad */
            {8'h00}, /* 0xc6ac */
            {8'h00}, /* 0xc6ab */
            {8'h00}, /* 0xc6aa */
            {8'h00}, /* 0xc6a9 */
            {8'h00}, /* 0xc6a8 */
            {8'h00}, /* 0xc6a7 */
            {8'h00}, /* 0xc6a6 */
            {8'h00}, /* 0xc6a5 */
            {8'h00}, /* 0xc6a4 */
            {8'h00}, /* 0xc6a3 */
            {8'h00}, /* 0xc6a2 */
            {8'h00}, /* 0xc6a1 */
            {8'h00}, /* 0xc6a0 */
            {8'h00}, /* 0xc69f */
            {8'h00}, /* 0xc69e */
            {8'h00}, /* 0xc69d */
            {8'h00}, /* 0xc69c */
            {8'h00}, /* 0xc69b */
            {8'h00}, /* 0xc69a */
            {8'h00}, /* 0xc699 */
            {8'h00}, /* 0xc698 */
            {8'h00}, /* 0xc697 */
            {8'h00}, /* 0xc696 */
            {8'h00}, /* 0xc695 */
            {8'h00}, /* 0xc694 */
            {8'h00}, /* 0xc693 */
            {8'h00}, /* 0xc692 */
            {8'h00}, /* 0xc691 */
            {8'h00}, /* 0xc690 */
            {8'h00}, /* 0xc68f */
            {8'h00}, /* 0xc68e */
            {8'h00}, /* 0xc68d */
            {8'h00}, /* 0xc68c */
            {8'h00}, /* 0xc68b */
            {8'h00}, /* 0xc68a */
            {8'h00}, /* 0xc689 */
            {8'h00}, /* 0xc688 */
            {8'h00}, /* 0xc687 */
            {8'h00}, /* 0xc686 */
            {8'h00}, /* 0xc685 */
            {8'h00}, /* 0xc684 */
            {8'h00}, /* 0xc683 */
            {8'h00}, /* 0xc682 */
            {8'h00}, /* 0xc681 */
            {8'h00}, /* 0xc680 */
            {8'h00}, /* 0xc67f */
            {8'h00}, /* 0xc67e */
            {8'h00}, /* 0xc67d */
            {8'h00}, /* 0xc67c */
            {8'h00}, /* 0xc67b */
            {8'h00}, /* 0xc67a */
            {8'h00}, /* 0xc679 */
            {8'h00}, /* 0xc678 */
            {8'h00}, /* 0xc677 */
            {8'h00}, /* 0xc676 */
            {8'h00}, /* 0xc675 */
            {8'h00}, /* 0xc674 */
            {8'h00}, /* 0xc673 */
            {8'h00}, /* 0xc672 */
            {8'h00}, /* 0xc671 */
            {8'h00}, /* 0xc670 */
            {8'h00}, /* 0xc66f */
            {8'h00}, /* 0xc66e */
            {8'h00}, /* 0xc66d */
            {8'h00}, /* 0xc66c */
            {8'h00}, /* 0xc66b */
            {8'h00}, /* 0xc66a */
            {8'h00}, /* 0xc669 */
            {8'h00}, /* 0xc668 */
            {8'h00}, /* 0xc667 */
            {8'h00}, /* 0xc666 */
            {8'h00}, /* 0xc665 */
            {8'h00}, /* 0xc664 */
            {8'h00}, /* 0xc663 */
            {8'h00}, /* 0xc662 */
            {8'h00}, /* 0xc661 */
            {8'h00}, /* 0xc660 */
            {8'h00}, /* 0xc65f */
            {8'h00}, /* 0xc65e */
            {8'h00}, /* 0xc65d */
            {8'h00}, /* 0xc65c */
            {8'h00}, /* 0xc65b */
            {8'h00}, /* 0xc65a */
            {8'h00}, /* 0xc659 */
            {8'h00}, /* 0xc658 */
            {8'h00}, /* 0xc657 */
            {8'h00}, /* 0xc656 */
            {8'h00}, /* 0xc655 */
            {8'h00}, /* 0xc654 */
            {8'h00}, /* 0xc653 */
            {8'h00}, /* 0xc652 */
            {8'h00}, /* 0xc651 */
            {8'h00}, /* 0xc650 */
            {8'h00}, /* 0xc64f */
            {8'h00}, /* 0xc64e */
            {8'h00}, /* 0xc64d */
            {8'h00}, /* 0xc64c */
            {8'h00}, /* 0xc64b */
            {8'h00}, /* 0xc64a */
            {8'h00}, /* 0xc649 */
            {8'h00}, /* 0xc648 */
            {8'h00}, /* 0xc647 */
            {8'h00}, /* 0xc646 */
            {8'h00}, /* 0xc645 */
            {8'h00}, /* 0xc644 */
            {8'h00}, /* 0xc643 */
            {8'h00}, /* 0xc642 */
            {8'h00}, /* 0xc641 */
            {8'h00}, /* 0xc640 */
            {8'h00}, /* 0xc63f */
            {8'h00}, /* 0xc63e */
            {8'h00}, /* 0xc63d */
            {8'h00}, /* 0xc63c */
            {8'h00}, /* 0xc63b */
            {8'h00}, /* 0xc63a */
            {8'h00}, /* 0xc639 */
            {8'h00}, /* 0xc638 */
            {8'h00}, /* 0xc637 */
            {8'h00}, /* 0xc636 */
            {8'h00}, /* 0xc635 */
            {8'h00}, /* 0xc634 */
            {8'h00}, /* 0xc633 */
            {8'h00}, /* 0xc632 */
            {8'h00}, /* 0xc631 */
            {8'h00}, /* 0xc630 */
            {8'h00}, /* 0xc62f */
            {8'h00}, /* 0xc62e */
            {8'h00}, /* 0xc62d */
            {8'h00}, /* 0xc62c */
            {8'h00}, /* 0xc62b */
            {8'h00}, /* 0xc62a */
            {8'h00}, /* 0xc629 */
            {8'h00}, /* 0xc628 */
            {8'h00}, /* 0xc627 */
            {8'h00}, /* 0xc626 */
            {8'h00}, /* 0xc625 */
            {8'h00}, /* 0xc624 */
            {8'h00}, /* 0xc623 */
            {8'h00}, /* 0xc622 */
            {8'h00}, /* 0xc621 */
            {8'h00}, /* 0xc620 */
            {8'h00}, /* 0xc61f */
            {8'h00}, /* 0xc61e */
            {8'h00}, /* 0xc61d */
            {8'h00}, /* 0xc61c */
            {8'h00}, /* 0xc61b */
            {8'h00}, /* 0xc61a */
            {8'h00}, /* 0xc619 */
            {8'h00}, /* 0xc618 */
            {8'h00}, /* 0xc617 */
            {8'h00}, /* 0xc616 */
            {8'h00}, /* 0xc615 */
            {8'h00}, /* 0xc614 */
            {8'h00}, /* 0xc613 */
            {8'h00}, /* 0xc612 */
            {8'h00}, /* 0xc611 */
            {8'h00}, /* 0xc610 */
            {8'h00}, /* 0xc60f */
            {8'h00}, /* 0xc60e */
            {8'h00}, /* 0xc60d */
            {8'h00}, /* 0xc60c */
            {8'h00}, /* 0xc60b */
            {8'h00}, /* 0xc60a */
            {8'h00}, /* 0xc609 */
            {8'h00}, /* 0xc608 */
            {8'h00}, /* 0xc607 */
            {8'h00}, /* 0xc606 */
            {8'h00}, /* 0xc605 */
            {8'h00}, /* 0xc604 */
            {8'h00}, /* 0xc603 */
            {8'h00}, /* 0xc602 */
            {8'h00}, /* 0xc601 */
            {8'h00}, /* 0xc600 */
            {8'h00}, /* 0xc5ff */
            {8'h00}, /* 0xc5fe */
            {8'h00}, /* 0xc5fd */
            {8'h00}, /* 0xc5fc */
            {8'h00}, /* 0xc5fb */
            {8'h00}, /* 0xc5fa */
            {8'h00}, /* 0xc5f9 */
            {8'h00}, /* 0xc5f8 */
            {8'h00}, /* 0xc5f7 */
            {8'h00}, /* 0xc5f6 */
            {8'h00}, /* 0xc5f5 */
            {8'h00}, /* 0xc5f4 */
            {8'h00}, /* 0xc5f3 */
            {8'h00}, /* 0xc5f2 */
            {8'h00}, /* 0xc5f1 */
            {8'h00}, /* 0xc5f0 */
            {8'h00}, /* 0xc5ef */
            {8'h00}, /* 0xc5ee */
            {8'h00}, /* 0xc5ed */
            {8'h00}, /* 0xc5ec */
            {8'h00}, /* 0xc5eb */
            {8'h00}, /* 0xc5ea */
            {8'h00}, /* 0xc5e9 */
            {8'h00}, /* 0xc5e8 */
            {8'h00}, /* 0xc5e7 */
            {8'h00}, /* 0xc5e6 */
            {8'h00}, /* 0xc5e5 */
            {8'h00}, /* 0xc5e4 */
            {8'h00}, /* 0xc5e3 */
            {8'h00}, /* 0xc5e2 */
            {8'h00}, /* 0xc5e1 */
            {8'h00}, /* 0xc5e0 */
            {8'h00}, /* 0xc5df */
            {8'h00}, /* 0xc5de */
            {8'h00}, /* 0xc5dd */
            {8'h00}, /* 0xc5dc */
            {8'h00}, /* 0xc5db */
            {8'h00}, /* 0xc5da */
            {8'h00}, /* 0xc5d9 */
            {8'h00}, /* 0xc5d8 */
            {8'h00}, /* 0xc5d7 */
            {8'h00}, /* 0xc5d6 */
            {8'h00}, /* 0xc5d5 */
            {8'h00}, /* 0xc5d4 */
            {8'h00}, /* 0xc5d3 */
            {8'h00}, /* 0xc5d2 */
            {8'h00}, /* 0xc5d1 */
            {8'h00}, /* 0xc5d0 */
            {8'h00}, /* 0xc5cf */
            {8'h00}, /* 0xc5ce */
            {8'h00}, /* 0xc5cd */
            {8'h00}, /* 0xc5cc */
            {8'h00}, /* 0xc5cb */
            {8'h00}, /* 0xc5ca */
            {8'h00}, /* 0xc5c9 */
            {8'h00}, /* 0xc5c8 */
            {8'h00}, /* 0xc5c7 */
            {8'h00}, /* 0xc5c6 */
            {8'h00}, /* 0xc5c5 */
            {8'h00}, /* 0xc5c4 */
            {8'h00}, /* 0xc5c3 */
            {8'h00}, /* 0xc5c2 */
            {8'h00}, /* 0xc5c1 */
            {8'h00}, /* 0xc5c0 */
            {8'h00}, /* 0xc5bf */
            {8'h00}, /* 0xc5be */
            {8'h00}, /* 0xc5bd */
            {8'h00}, /* 0xc5bc */
            {8'h00}, /* 0xc5bb */
            {8'h00}, /* 0xc5ba */
            {8'h00}, /* 0xc5b9 */
            {8'h00}, /* 0xc5b8 */
            {8'h00}, /* 0xc5b7 */
            {8'h00}, /* 0xc5b6 */
            {8'h00}, /* 0xc5b5 */
            {8'h00}, /* 0xc5b4 */
            {8'h00}, /* 0xc5b3 */
            {8'h00}, /* 0xc5b2 */
            {8'h00}, /* 0xc5b1 */
            {8'h00}, /* 0xc5b0 */
            {8'h00}, /* 0xc5af */
            {8'h00}, /* 0xc5ae */
            {8'h00}, /* 0xc5ad */
            {8'h00}, /* 0xc5ac */
            {8'h00}, /* 0xc5ab */
            {8'h00}, /* 0xc5aa */
            {8'h00}, /* 0xc5a9 */
            {8'h00}, /* 0xc5a8 */
            {8'h00}, /* 0xc5a7 */
            {8'h00}, /* 0xc5a6 */
            {8'h00}, /* 0xc5a5 */
            {8'h00}, /* 0xc5a4 */
            {8'h00}, /* 0xc5a3 */
            {8'h00}, /* 0xc5a2 */
            {8'h00}, /* 0xc5a1 */
            {8'h00}, /* 0xc5a0 */
            {8'h00}, /* 0xc59f */
            {8'h00}, /* 0xc59e */
            {8'h00}, /* 0xc59d */
            {8'h00}, /* 0xc59c */
            {8'h00}, /* 0xc59b */
            {8'h00}, /* 0xc59a */
            {8'h00}, /* 0xc599 */
            {8'h00}, /* 0xc598 */
            {8'h00}, /* 0xc597 */
            {8'h00}, /* 0xc596 */
            {8'h00}, /* 0xc595 */
            {8'h00}, /* 0xc594 */
            {8'h00}, /* 0xc593 */
            {8'h00}, /* 0xc592 */
            {8'h00}, /* 0xc591 */
            {8'h00}, /* 0xc590 */
            {8'h00}, /* 0xc58f */
            {8'h00}, /* 0xc58e */
            {8'h00}, /* 0xc58d */
            {8'h00}, /* 0xc58c */
            {8'h00}, /* 0xc58b */
            {8'h00}, /* 0xc58a */
            {8'h00}, /* 0xc589 */
            {8'h00}, /* 0xc588 */
            {8'h00}, /* 0xc587 */
            {8'h00}, /* 0xc586 */
            {8'h00}, /* 0xc585 */
            {8'h00}, /* 0xc584 */
            {8'h00}, /* 0xc583 */
            {8'h00}, /* 0xc582 */
            {8'h00}, /* 0xc581 */
            {8'h00}, /* 0xc580 */
            {8'h00}, /* 0xc57f */
            {8'h00}, /* 0xc57e */
            {8'h00}, /* 0xc57d */
            {8'h00}, /* 0xc57c */
            {8'h00}, /* 0xc57b */
            {8'h00}, /* 0xc57a */
            {8'h00}, /* 0xc579 */
            {8'h00}, /* 0xc578 */
            {8'h00}, /* 0xc577 */
            {8'h00}, /* 0xc576 */
            {8'h00}, /* 0xc575 */
            {8'h00}, /* 0xc574 */
            {8'h00}, /* 0xc573 */
            {8'h00}, /* 0xc572 */
            {8'h00}, /* 0xc571 */
            {8'h00}, /* 0xc570 */
            {8'h00}, /* 0xc56f */
            {8'h00}, /* 0xc56e */
            {8'h00}, /* 0xc56d */
            {8'h00}, /* 0xc56c */
            {8'h00}, /* 0xc56b */
            {8'h00}, /* 0xc56a */
            {8'h00}, /* 0xc569 */
            {8'h00}, /* 0xc568 */
            {8'h00}, /* 0xc567 */
            {8'h00}, /* 0xc566 */
            {8'h00}, /* 0xc565 */
            {8'h00}, /* 0xc564 */
            {8'h00}, /* 0xc563 */
            {8'h00}, /* 0xc562 */
            {8'h00}, /* 0xc561 */
            {8'h00}, /* 0xc560 */
            {8'h00}, /* 0xc55f */
            {8'h00}, /* 0xc55e */
            {8'h00}, /* 0xc55d */
            {8'h00}, /* 0xc55c */
            {8'h00}, /* 0xc55b */
            {8'h00}, /* 0xc55a */
            {8'h00}, /* 0xc559 */
            {8'h00}, /* 0xc558 */
            {8'h00}, /* 0xc557 */
            {8'h00}, /* 0xc556 */
            {8'h00}, /* 0xc555 */
            {8'h00}, /* 0xc554 */
            {8'h00}, /* 0xc553 */
            {8'h00}, /* 0xc552 */
            {8'h00}, /* 0xc551 */
            {8'h00}, /* 0xc550 */
            {8'h00}, /* 0xc54f */
            {8'h00}, /* 0xc54e */
            {8'h00}, /* 0xc54d */
            {8'h00}, /* 0xc54c */
            {8'h00}, /* 0xc54b */
            {8'h00}, /* 0xc54a */
            {8'h00}, /* 0xc549 */
            {8'h00}, /* 0xc548 */
            {8'h00}, /* 0xc547 */
            {8'h00}, /* 0xc546 */
            {8'h00}, /* 0xc545 */
            {8'h00}, /* 0xc544 */
            {8'h00}, /* 0xc543 */
            {8'h00}, /* 0xc542 */
            {8'h00}, /* 0xc541 */
            {8'h00}, /* 0xc540 */
            {8'h00}, /* 0xc53f */
            {8'h00}, /* 0xc53e */
            {8'h00}, /* 0xc53d */
            {8'h00}, /* 0xc53c */
            {8'h00}, /* 0xc53b */
            {8'h00}, /* 0xc53a */
            {8'h00}, /* 0xc539 */
            {8'h00}, /* 0xc538 */
            {8'h00}, /* 0xc537 */
            {8'h00}, /* 0xc536 */
            {8'h00}, /* 0xc535 */
            {8'h00}, /* 0xc534 */
            {8'h00}, /* 0xc533 */
            {8'h00}, /* 0xc532 */
            {8'h00}, /* 0xc531 */
            {8'h00}, /* 0xc530 */
            {8'h00}, /* 0xc52f */
            {8'h00}, /* 0xc52e */
            {8'h00}, /* 0xc52d */
            {8'h00}, /* 0xc52c */
            {8'h00}, /* 0xc52b */
            {8'h00}, /* 0xc52a */
            {8'h00}, /* 0xc529 */
            {8'h00}, /* 0xc528 */
            {8'h00}, /* 0xc527 */
            {8'h00}, /* 0xc526 */
            {8'h00}, /* 0xc525 */
            {8'h00}, /* 0xc524 */
            {8'h00}, /* 0xc523 */
            {8'h00}, /* 0xc522 */
            {8'h00}, /* 0xc521 */
            {8'h00}, /* 0xc520 */
            {8'h00}, /* 0xc51f */
            {8'h00}, /* 0xc51e */
            {8'h00}, /* 0xc51d */
            {8'h00}, /* 0xc51c */
            {8'h00}, /* 0xc51b */
            {8'h00}, /* 0xc51a */
            {8'h00}, /* 0xc519 */
            {8'h00}, /* 0xc518 */
            {8'h00}, /* 0xc517 */
            {8'h00}, /* 0xc516 */
            {8'h00}, /* 0xc515 */
            {8'h00}, /* 0xc514 */
            {8'h00}, /* 0xc513 */
            {8'h00}, /* 0xc512 */
            {8'h00}, /* 0xc511 */
            {8'h00}, /* 0xc510 */
            {8'h00}, /* 0xc50f */
            {8'h00}, /* 0xc50e */
            {8'h00}, /* 0xc50d */
            {8'h00}, /* 0xc50c */
            {8'h00}, /* 0xc50b */
            {8'h00}, /* 0xc50a */
            {8'h00}, /* 0xc509 */
            {8'h00}, /* 0xc508 */
            {8'h00}, /* 0xc507 */
            {8'h00}, /* 0xc506 */
            {8'h00}, /* 0xc505 */
            {8'h00}, /* 0xc504 */
            {8'h00}, /* 0xc503 */
            {8'h00}, /* 0xc502 */
            {8'h00}, /* 0xc501 */
            {8'h00}, /* 0xc500 */
            {8'h00}, /* 0xc4ff */
            {8'h00}, /* 0xc4fe */
            {8'h00}, /* 0xc4fd */
            {8'h00}, /* 0xc4fc */
            {8'h00}, /* 0xc4fb */
            {8'h00}, /* 0xc4fa */
            {8'h00}, /* 0xc4f9 */
            {8'h00}, /* 0xc4f8 */
            {8'h00}, /* 0xc4f7 */
            {8'h00}, /* 0xc4f6 */
            {8'h00}, /* 0xc4f5 */
            {8'h00}, /* 0xc4f4 */
            {8'h00}, /* 0xc4f3 */
            {8'h00}, /* 0xc4f2 */
            {8'h00}, /* 0xc4f1 */
            {8'h00}, /* 0xc4f0 */
            {8'h00}, /* 0xc4ef */
            {8'h00}, /* 0xc4ee */
            {8'h00}, /* 0xc4ed */
            {8'h00}, /* 0xc4ec */
            {8'h00}, /* 0xc4eb */
            {8'h00}, /* 0xc4ea */
            {8'h00}, /* 0xc4e9 */
            {8'h00}, /* 0xc4e8 */
            {8'h00}, /* 0xc4e7 */
            {8'h00}, /* 0xc4e6 */
            {8'h00}, /* 0xc4e5 */
            {8'h00}, /* 0xc4e4 */
            {8'h00}, /* 0xc4e3 */
            {8'h00}, /* 0xc4e2 */
            {8'h00}, /* 0xc4e1 */
            {8'h00}, /* 0xc4e0 */
            {8'h00}, /* 0xc4df */
            {8'h00}, /* 0xc4de */
            {8'h00}, /* 0xc4dd */
            {8'h00}, /* 0xc4dc */
            {8'h00}, /* 0xc4db */
            {8'h00}, /* 0xc4da */
            {8'h00}, /* 0xc4d9 */
            {8'h00}, /* 0xc4d8 */
            {8'h00}, /* 0xc4d7 */
            {8'h00}, /* 0xc4d6 */
            {8'h00}, /* 0xc4d5 */
            {8'h00}, /* 0xc4d4 */
            {8'h00}, /* 0xc4d3 */
            {8'h00}, /* 0xc4d2 */
            {8'h00}, /* 0xc4d1 */
            {8'h00}, /* 0xc4d0 */
            {8'h00}, /* 0xc4cf */
            {8'h00}, /* 0xc4ce */
            {8'h00}, /* 0xc4cd */
            {8'h00}, /* 0xc4cc */
            {8'h00}, /* 0xc4cb */
            {8'h00}, /* 0xc4ca */
            {8'h00}, /* 0xc4c9 */
            {8'h00}, /* 0xc4c8 */
            {8'h00}, /* 0xc4c7 */
            {8'h00}, /* 0xc4c6 */
            {8'h00}, /* 0xc4c5 */
            {8'h00}, /* 0xc4c4 */
            {8'h00}, /* 0xc4c3 */
            {8'h00}, /* 0xc4c2 */
            {8'h00}, /* 0xc4c1 */
            {8'h00}, /* 0xc4c0 */
            {8'h00}, /* 0xc4bf */
            {8'h00}, /* 0xc4be */
            {8'h00}, /* 0xc4bd */
            {8'h00}, /* 0xc4bc */
            {8'h00}, /* 0xc4bb */
            {8'h00}, /* 0xc4ba */
            {8'h00}, /* 0xc4b9 */
            {8'h00}, /* 0xc4b8 */
            {8'h00}, /* 0xc4b7 */
            {8'h00}, /* 0xc4b6 */
            {8'h00}, /* 0xc4b5 */
            {8'h00}, /* 0xc4b4 */
            {8'h00}, /* 0xc4b3 */
            {8'h00}, /* 0xc4b2 */
            {8'h00}, /* 0xc4b1 */
            {8'h00}, /* 0xc4b0 */
            {8'h00}, /* 0xc4af */
            {8'h00}, /* 0xc4ae */
            {8'h00}, /* 0xc4ad */
            {8'h00}, /* 0xc4ac */
            {8'h00}, /* 0xc4ab */
            {8'h00}, /* 0xc4aa */
            {8'h00}, /* 0xc4a9 */
            {8'h00}, /* 0xc4a8 */
            {8'h00}, /* 0xc4a7 */
            {8'h00}, /* 0xc4a6 */
            {8'h00}, /* 0xc4a5 */
            {8'h00}, /* 0xc4a4 */
            {8'h00}, /* 0xc4a3 */
            {8'h00}, /* 0xc4a2 */
            {8'h00}, /* 0xc4a1 */
            {8'h00}, /* 0xc4a0 */
            {8'h00}, /* 0xc49f */
            {8'h00}, /* 0xc49e */
            {8'h00}, /* 0xc49d */
            {8'h00}, /* 0xc49c */
            {8'h00}, /* 0xc49b */
            {8'h00}, /* 0xc49a */
            {8'h00}, /* 0xc499 */
            {8'h00}, /* 0xc498 */
            {8'h00}, /* 0xc497 */
            {8'h00}, /* 0xc496 */
            {8'h00}, /* 0xc495 */
            {8'h00}, /* 0xc494 */
            {8'h00}, /* 0xc493 */
            {8'h00}, /* 0xc492 */
            {8'h00}, /* 0xc491 */
            {8'h00}, /* 0xc490 */
            {8'h00}, /* 0xc48f */
            {8'h00}, /* 0xc48e */
            {8'h00}, /* 0xc48d */
            {8'h00}, /* 0xc48c */
            {8'h00}, /* 0xc48b */
            {8'h00}, /* 0xc48a */
            {8'h00}, /* 0xc489 */
            {8'h00}, /* 0xc488 */
            {8'h00}, /* 0xc487 */
            {8'h00}, /* 0xc486 */
            {8'h00}, /* 0xc485 */
            {8'h00}, /* 0xc484 */
            {8'h00}, /* 0xc483 */
            {8'h00}, /* 0xc482 */
            {8'h00}, /* 0xc481 */
            {8'h00}, /* 0xc480 */
            {8'h00}, /* 0xc47f */
            {8'h00}, /* 0xc47e */
            {8'h00}, /* 0xc47d */
            {8'h00}, /* 0xc47c */
            {8'h00}, /* 0xc47b */
            {8'h00}, /* 0xc47a */
            {8'h00}, /* 0xc479 */
            {8'h00}, /* 0xc478 */
            {8'h00}, /* 0xc477 */
            {8'h00}, /* 0xc476 */
            {8'h00}, /* 0xc475 */
            {8'h00}, /* 0xc474 */
            {8'h00}, /* 0xc473 */
            {8'h00}, /* 0xc472 */
            {8'h00}, /* 0xc471 */
            {8'h00}, /* 0xc470 */
            {8'h00}, /* 0xc46f */
            {8'h00}, /* 0xc46e */
            {8'h00}, /* 0xc46d */
            {8'h00}, /* 0xc46c */
            {8'h00}, /* 0xc46b */
            {8'h00}, /* 0xc46a */
            {8'h00}, /* 0xc469 */
            {8'h00}, /* 0xc468 */
            {8'h00}, /* 0xc467 */
            {8'h00}, /* 0xc466 */
            {8'h00}, /* 0xc465 */
            {8'h00}, /* 0xc464 */
            {8'h00}, /* 0xc463 */
            {8'h00}, /* 0xc462 */
            {8'h00}, /* 0xc461 */
            {8'h00}, /* 0xc460 */
            {8'h00}, /* 0xc45f */
            {8'h00}, /* 0xc45e */
            {8'h00}, /* 0xc45d */
            {8'h00}, /* 0xc45c */
            {8'h00}, /* 0xc45b */
            {8'h00}, /* 0xc45a */
            {8'h00}, /* 0xc459 */
            {8'h00}, /* 0xc458 */
            {8'h00}, /* 0xc457 */
            {8'h00}, /* 0xc456 */
            {8'h00}, /* 0xc455 */
            {8'h00}, /* 0xc454 */
            {8'h00}, /* 0xc453 */
            {8'h00}, /* 0xc452 */
            {8'h00}, /* 0xc451 */
            {8'h00}, /* 0xc450 */
            {8'h00}, /* 0xc44f */
            {8'h00}, /* 0xc44e */
            {8'h00}, /* 0xc44d */
            {8'h00}, /* 0xc44c */
            {8'h00}, /* 0xc44b */
            {8'h00}, /* 0xc44a */
            {8'h00}, /* 0xc449 */
            {8'h00}, /* 0xc448 */
            {8'h00}, /* 0xc447 */
            {8'h00}, /* 0xc446 */
            {8'h00}, /* 0xc445 */
            {8'h00}, /* 0xc444 */
            {8'h00}, /* 0xc443 */
            {8'h00}, /* 0xc442 */
            {8'h00}, /* 0xc441 */
            {8'h00}, /* 0xc440 */
            {8'h00}, /* 0xc43f */
            {8'h00}, /* 0xc43e */
            {8'h00}, /* 0xc43d */
            {8'h00}, /* 0xc43c */
            {8'h00}, /* 0xc43b */
            {8'h00}, /* 0xc43a */
            {8'h00}, /* 0xc439 */
            {8'h00}, /* 0xc438 */
            {8'h00}, /* 0xc437 */
            {8'h00}, /* 0xc436 */
            {8'h00}, /* 0xc435 */
            {8'h00}, /* 0xc434 */
            {8'h00}, /* 0xc433 */
            {8'h00}, /* 0xc432 */
            {8'h00}, /* 0xc431 */
            {8'h00}, /* 0xc430 */
            {8'h00}, /* 0xc42f */
            {8'h00}, /* 0xc42e */
            {8'h00}, /* 0xc42d */
            {8'h00}, /* 0xc42c */
            {8'h00}, /* 0xc42b */
            {8'h00}, /* 0xc42a */
            {8'h00}, /* 0xc429 */
            {8'h00}, /* 0xc428 */
            {8'h00}, /* 0xc427 */
            {8'h00}, /* 0xc426 */
            {8'h00}, /* 0xc425 */
            {8'h00}, /* 0xc424 */
            {8'h00}, /* 0xc423 */
            {8'h00}, /* 0xc422 */
            {8'h00}, /* 0xc421 */
            {8'h00}, /* 0xc420 */
            {8'h00}, /* 0xc41f */
            {8'h00}, /* 0xc41e */
            {8'h00}, /* 0xc41d */
            {8'h00}, /* 0xc41c */
            {8'h00}, /* 0xc41b */
            {8'h00}, /* 0xc41a */
            {8'h00}, /* 0xc419 */
            {8'h00}, /* 0xc418 */
            {8'h00}, /* 0xc417 */
            {8'h00}, /* 0xc416 */
            {8'h00}, /* 0xc415 */
            {8'h00}, /* 0xc414 */
            {8'h00}, /* 0xc413 */
            {8'h00}, /* 0xc412 */
            {8'h00}, /* 0xc411 */
            {8'h00}, /* 0xc410 */
            {8'h00}, /* 0xc40f */
            {8'h00}, /* 0xc40e */
            {8'h00}, /* 0xc40d */
            {8'h00}, /* 0xc40c */
            {8'h00}, /* 0xc40b */
            {8'h00}, /* 0xc40a */
            {8'h00}, /* 0xc409 */
            {8'h00}, /* 0xc408 */
            {8'h00}, /* 0xc407 */
            {8'h00}, /* 0xc406 */
            {8'h00}, /* 0xc405 */
            {8'h00}, /* 0xc404 */
            {8'h00}, /* 0xc403 */
            {8'h00}, /* 0xc402 */
            {8'h00}, /* 0xc401 */
            {8'h00}, /* 0xc400 */
            {8'h00}, /* 0xc3ff */
            {8'h00}, /* 0xc3fe */
            {8'h00}, /* 0xc3fd */
            {8'h00}, /* 0xc3fc */
            {8'h00}, /* 0xc3fb */
            {8'h00}, /* 0xc3fa */
            {8'h00}, /* 0xc3f9 */
            {8'h00}, /* 0xc3f8 */
            {8'h00}, /* 0xc3f7 */
            {8'h00}, /* 0xc3f6 */
            {8'h00}, /* 0xc3f5 */
            {8'h00}, /* 0xc3f4 */
            {8'h00}, /* 0xc3f3 */
            {8'h00}, /* 0xc3f2 */
            {8'h00}, /* 0xc3f1 */
            {8'h00}, /* 0xc3f0 */
            {8'h00}, /* 0xc3ef */
            {8'h00}, /* 0xc3ee */
            {8'h00}, /* 0xc3ed */
            {8'h00}, /* 0xc3ec */
            {8'h00}, /* 0xc3eb */
            {8'h00}, /* 0xc3ea */
            {8'h00}, /* 0xc3e9 */
            {8'h00}, /* 0xc3e8 */
            {8'h00}, /* 0xc3e7 */
            {8'h00}, /* 0xc3e6 */
            {8'h00}, /* 0xc3e5 */
            {8'h00}, /* 0xc3e4 */
            {8'h00}, /* 0xc3e3 */
            {8'h00}, /* 0xc3e2 */
            {8'h00}, /* 0xc3e1 */
            {8'h00}, /* 0xc3e0 */
            {8'h00}, /* 0xc3df */
            {8'h00}, /* 0xc3de */
            {8'h00}, /* 0xc3dd */
            {8'h00}, /* 0xc3dc */
            {8'h00}, /* 0xc3db */
            {8'h00}, /* 0xc3da */
            {8'h00}, /* 0xc3d9 */
            {8'h00}, /* 0xc3d8 */
            {8'h00}, /* 0xc3d7 */
            {8'h00}, /* 0xc3d6 */
            {8'h00}, /* 0xc3d5 */
            {8'h00}, /* 0xc3d4 */
            {8'h00}, /* 0xc3d3 */
            {8'h00}, /* 0xc3d2 */
            {8'h00}, /* 0xc3d1 */
            {8'h00}, /* 0xc3d0 */
            {8'h00}, /* 0xc3cf */
            {8'h00}, /* 0xc3ce */
            {8'h00}, /* 0xc3cd */
            {8'h00}, /* 0xc3cc */
            {8'h00}, /* 0xc3cb */
            {8'h00}, /* 0xc3ca */
            {8'h00}, /* 0xc3c9 */
            {8'h00}, /* 0xc3c8 */
            {8'h00}, /* 0xc3c7 */
            {8'h00}, /* 0xc3c6 */
            {8'h00}, /* 0xc3c5 */
            {8'h00}, /* 0xc3c4 */
            {8'h00}, /* 0xc3c3 */
            {8'h00}, /* 0xc3c2 */
            {8'h00}, /* 0xc3c1 */
            {8'h00}, /* 0xc3c0 */
            {8'h00}, /* 0xc3bf */
            {8'h00}, /* 0xc3be */
            {8'h00}, /* 0xc3bd */
            {8'h00}, /* 0xc3bc */
            {8'h00}, /* 0xc3bb */
            {8'h00}, /* 0xc3ba */
            {8'h00}, /* 0xc3b9 */
            {8'h00}, /* 0xc3b8 */
            {8'h00}, /* 0xc3b7 */
            {8'h00}, /* 0xc3b6 */
            {8'h00}, /* 0xc3b5 */
            {8'h00}, /* 0xc3b4 */
            {8'h00}, /* 0xc3b3 */
            {8'h00}, /* 0xc3b2 */
            {8'h00}, /* 0xc3b1 */
            {8'h00}, /* 0xc3b0 */
            {8'h00}, /* 0xc3af */
            {8'h00}, /* 0xc3ae */
            {8'h00}, /* 0xc3ad */
            {8'h00}, /* 0xc3ac */
            {8'h00}, /* 0xc3ab */
            {8'h00}, /* 0xc3aa */
            {8'h00}, /* 0xc3a9 */
            {8'h00}, /* 0xc3a8 */
            {8'h00}, /* 0xc3a7 */
            {8'h00}, /* 0xc3a6 */
            {8'h00}, /* 0xc3a5 */
            {8'h00}, /* 0xc3a4 */
            {8'h00}, /* 0xc3a3 */
            {8'h00}, /* 0xc3a2 */
            {8'h00}, /* 0xc3a1 */
            {8'h00}, /* 0xc3a0 */
            {8'h00}, /* 0xc39f */
            {8'h00}, /* 0xc39e */
            {8'h00}, /* 0xc39d */
            {8'h00}, /* 0xc39c */
            {8'h00}, /* 0xc39b */
            {8'h00}, /* 0xc39a */
            {8'h00}, /* 0xc399 */
            {8'h00}, /* 0xc398 */
            {8'h00}, /* 0xc397 */
            {8'h00}, /* 0xc396 */
            {8'h00}, /* 0xc395 */
            {8'h00}, /* 0xc394 */
            {8'h00}, /* 0xc393 */
            {8'h00}, /* 0xc392 */
            {8'h00}, /* 0xc391 */
            {8'h00}, /* 0xc390 */
            {8'h00}, /* 0xc38f */
            {8'h00}, /* 0xc38e */
            {8'h00}, /* 0xc38d */
            {8'h00}, /* 0xc38c */
            {8'h00}, /* 0xc38b */
            {8'h00}, /* 0xc38a */
            {8'h00}, /* 0xc389 */
            {8'h00}, /* 0xc388 */
            {8'h00}, /* 0xc387 */
            {8'h00}, /* 0xc386 */
            {8'h00}, /* 0xc385 */
            {8'h00}, /* 0xc384 */
            {8'h00}, /* 0xc383 */
            {8'h00}, /* 0xc382 */
            {8'h00}, /* 0xc381 */
            {8'h00}, /* 0xc380 */
            {8'h00}, /* 0xc37f */
            {8'h00}, /* 0xc37e */
            {8'h00}, /* 0xc37d */
            {8'h00}, /* 0xc37c */
            {8'h00}, /* 0xc37b */
            {8'h00}, /* 0xc37a */
            {8'h00}, /* 0xc379 */
            {8'h00}, /* 0xc378 */
            {8'h00}, /* 0xc377 */
            {8'h00}, /* 0xc376 */
            {8'h00}, /* 0xc375 */
            {8'h00}, /* 0xc374 */
            {8'h00}, /* 0xc373 */
            {8'h00}, /* 0xc372 */
            {8'h00}, /* 0xc371 */
            {8'h00}, /* 0xc370 */
            {8'h00}, /* 0xc36f */
            {8'h00}, /* 0xc36e */
            {8'h00}, /* 0xc36d */
            {8'h00}, /* 0xc36c */
            {8'h00}, /* 0xc36b */
            {8'h00}, /* 0xc36a */
            {8'h00}, /* 0xc369 */
            {8'h00}, /* 0xc368 */
            {8'h00}, /* 0xc367 */
            {8'h00}, /* 0xc366 */
            {8'h00}, /* 0xc365 */
            {8'h00}, /* 0xc364 */
            {8'h00}, /* 0xc363 */
            {8'h00}, /* 0xc362 */
            {8'h00}, /* 0xc361 */
            {8'h00}, /* 0xc360 */
            {8'h00}, /* 0xc35f */
            {8'h00}, /* 0xc35e */
            {8'h00}, /* 0xc35d */
            {8'h00}, /* 0xc35c */
            {8'h00}, /* 0xc35b */
            {8'h00}, /* 0xc35a */
            {8'h00}, /* 0xc359 */
            {8'h00}, /* 0xc358 */
            {8'h00}, /* 0xc357 */
            {8'h00}, /* 0xc356 */
            {8'h00}, /* 0xc355 */
            {8'h00}, /* 0xc354 */
            {8'h00}, /* 0xc353 */
            {8'h00}, /* 0xc352 */
            {8'h00}, /* 0xc351 */
            {8'h00}, /* 0xc350 */
            {8'h00}, /* 0xc34f */
            {8'h00}, /* 0xc34e */
            {8'h00}, /* 0xc34d */
            {8'h00}, /* 0xc34c */
            {8'h00}, /* 0xc34b */
            {8'h00}, /* 0xc34a */
            {8'h00}, /* 0xc349 */
            {8'h00}, /* 0xc348 */
            {8'h00}, /* 0xc347 */
            {8'h00}, /* 0xc346 */
            {8'h00}, /* 0xc345 */
            {8'h00}, /* 0xc344 */
            {8'h00}, /* 0xc343 */
            {8'h00}, /* 0xc342 */
            {8'h00}, /* 0xc341 */
            {8'h00}, /* 0xc340 */
            {8'h00}, /* 0xc33f */
            {8'h00}, /* 0xc33e */
            {8'h00}, /* 0xc33d */
            {8'h00}, /* 0xc33c */
            {8'h00}, /* 0xc33b */
            {8'h00}, /* 0xc33a */
            {8'h00}, /* 0xc339 */
            {8'h00}, /* 0xc338 */
            {8'h00}, /* 0xc337 */
            {8'h00}, /* 0xc336 */
            {8'h00}, /* 0xc335 */
            {8'h00}, /* 0xc334 */
            {8'h00}, /* 0xc333 */
            {8'h00}, /* 0xc332 */
            {8'h00}, /* 0xc331 */
            {8'h00}, /* 0xc330 */
            {8'h00}, /* 0xc32f */
            {8'h00}, /* 0xc32e */
            {8'h00}, /* 0xc32d */
            {8'h00}, /* 0xc32c */
            {8'h00}, /* 0xc32b */
            {8'h00}, /* 0xc32a */
            {8'h00}, /* 0xc329 */
            {8'h00}, /* 0xc328 */
            {8'h00}, /* 0xc327 */
            {8'h00}, /* 0xc326 */
            {8'h00}, /* 0xc325 */
            {8'h00}, /* 0xc324 */
            {8'h00}, /* 0xc323 */
            {8'h00}, /* 0xc322 */
            {8'h00}, /* 0xc321 */
            {8'h00}, /* 0xc320 */
            {8'h00}, /* 0xc31f */
            {8'h00}, /* 0xc31e */
            {8'h00}, /* 0xc31d */
            {8'h00}, /* 0xc31c */
            {8'h00}, /* 0xc31b */
            {8'h00}, /* 0xc31a */
            {8'h00}, /* 0xc319 */
            {8'h00}, /* 0xc318 */
            {8'h00}, /* 0xc317 */
            {8'h00}, /* 0xc316 */
            {8'h00}, /* 0xc315 */
            {8'h00}, /* 0xc314 */
            {8'h00}, /* 0xc313 */
            {8'h00}, /* 0xc312 */
            {8'h00}, /* 0xc311 */
            {8'h00}, /* 0xc310 */
            {8'h00}, /* 0xc30f */
            {8'h00}, /* 0xc30e */
            {8'h00}, /* 0xc30d */
            {8'h00}, /* 0xc30c */
            {8'h00}, /* 0xc30b */
            {8'h00}, /* 0xc30a */
            {8'h00}, /* 0xc309 */
            {8'h00}, /* 0xc308 */
            {8'h00}, /* 0xc307 */
            {8'h00}, /* 0xc306 */
            {8'h00}, /* 0xc305 */
            {8'h00}, /* 0xc304 */
            {8'h00}, /* 0xc303 */
            {8'h00}, /* 0xc302 */
            {8'h00}, /* 0xc301 */
            {8'h00}, /* 0xc300 */
            {8'h00}, /* 0xc2ff */
            {8'h00}, /* 0xc2fe */
            {8'h00}, /* 0xc2fd */
            {8'h00}, /* 0xc2fc */
            {8'h00}, /* 0xc2fb */
            {8'h00}, /* 0xc2fa */
            {8'h00}, /* 0xc2f9 */
            {8'h00}, /* 0xc2f8 */
            {8'h00}, /* 0xc2f7 */
            {8'h00}, /* 0xc2f6 */
            {8'h00}, /* 0xc2f5 */
            {8'h00}, /* 0xc2f4 */
            {8'h00}, /* 0xc2f3 */
            {8'h00}, /* 0xc2f2 */
            {8'h00}, /* 0xc2f1 */
            {8'h00}, /* 0xc2f0 */
            {8'h00}, /* 0xc2ef */
            {8'h00}, /* 0xc2ee */
            {8'h00}, /* 0xc2ed */
            {8'h00}, /* 0xc2ec */
            {8'h00}, /* 0xc2eb */
            {8'h00}, /* 0xc2ea */
            {8'h00}, /* 0xc2e9 */
            {8'h00}, /* 0xc2e8 */
            {8'h00}, /* 0xc2e7 */
            {8'h00}, /* 0xc2e6 */
            {8'h00}, /* 0xc2e5 */
            {8'h00}, /* 0xc2e4 */
            {8'h00}, /* 0xc2e3 */
            {8'h00}, /* 0xc2e2 */
            {8'h00}, /* 0xc2e1 */
            {8'h00}, /* 0xc2e0 */
            {8'h00}, /* 0xc2df */
            {8'h00}, /* 0xc2de */
            {8'h00}, /* 0xc2dd */
            {8'h00}, /* 0xc2dc */
            {8'h00}, /* 0xc2db */
            {8'h00}, /* 0xc2da */
            {8'h00}, /* 0xc2d9 */
            {8'h00}, /* 0xc2d8 */
            {8'h00}, /* 0xc2d7 */
            {8'h00}, /* 0xc2d6 */
            {8'h00}, /* 0xc2d5 */
            {8'h00}, /* 0xc2d4 */
            {8'h00}, /* 0xc2d3 */
            {8'h00}, /* 0xc2d2 */
            {8'h00}, /* 0xc2d1 */
            {8'h00}, /* 0xc2d0 */
            {8'h00}, /* 0xc2cf */
            {8'h00}, /* 0xc2ce */
            {8'h00}, /* 0xc2cd */
            {8'h00}, /* 0xc2cc */
            {8'h00}, /* 0xc2cb */
            {8'h00}, /* 0xc2ca */
            {8'h00}, /* 0xc2c9 */
            {8'h00}, /* 0xc2c8 */
            {8'h00}, /* 0xc2c7 */
            {8'h00}, /* 0xc2c6 */
            {8'h00}, /* 0xc2c5 */
            {8'h00}, /* 0xc2c4 */
            {8'h00}, /* 0xc2c3 */
            {8'h00}, /* 0xc2c2 */
            {8'h00}, /* 0xc2c1 */
            {8'h00}, /* 0xc2c0 */
            {8'h00}, /* 0xc2bf */
            {8'h00}, /* 0xc2be */
            {8'h00}, /* 0xc2bd */
            {8'h00}, /* 0xc2bc */
            {8'h00}, /* 0xc2bb */
            {8'h00}, /* 0xc2ba */
            {8'h00}, /* 0xc2b9 */
            {8'h00}, /* 0xc2b8 */
            {8'h00}, /* 0xc2b7 */
            {8'h00}, /* 0xc2b6 */
            {8'h00}, /* 0xc2b5 */
            {8'h00}, /* 0xc2b4 */
            {8'h00}, /* 0xc2b3 */
            {8'h00}, /* 0xc2b2 */
            {8'h00}, /* 0xc2b1 */
            {8'h00}, /* 0xc2b0 */
            {8'h00}, /* 0xc2af */
            {8'h00}, /* 0xc2ae */
            {8'h00}, /* 0xc2ad */
            {8'h00}, /* 0xc2ac */
            {8'h00}, /* 0xc2ab */
            {8'h00}, /* 0xc2aa */
            {8'h00}, /* 0xc2a9 */
            {8'h00}, /* 0xc2a8 */
            {8'h00}, /* 0xc2a7 */
            {8'h00}, /* 0xc2a6 */
            {8'h00}, /* 0xc2a5 */
            {8'h00}, /* 0xc2a4 */
            {8'h00}, /* 0xc2a3 */
            {8'h00}, /* 0xc2a2 */
            {8'h00}, /* 0xc2a1 */
            {8'h00}, /* 0xc2a0 */
            {8'h00}, /* 0xc29f */
            {8'h00}, /* 0xc29e */
            {8'h00}, /* 0xc29d */
            {8'h00}, /* 0xc29c */
            {8'h00}, /* 0xc29b */
            {8'h00}, /* 0xc29a */
            {8'h00}, /* 0xc299 */
            {8'h00}, /* 0xc298 */
            {8'h00}, /* 0xc297 */
            {8'h00}, /* 0xc296 */
            {8'h00}, /* 0xc295 */
            {8'h00}, /* 0xc294 */
            {8'h00}, /* 0xc293 */
            {8'h00}, /* 0xc292 */
            {8'h00}, /* 0xc291 */
            {8'h00}, /* 0xc290 */
            {8'h00}, /* 0xc28f */
            {8'h00}, /* 0xc28e */
            {8'h00}, /* 0xc28d */
            {8'h00}, /* 0xc28c */
            {8'h00}, /* 0xc28b */
            {8'h00}, /* 0xc28a */
            {8'h00}, /* 0xc289 */
            {8'h00}, /* 0xc288 */
            {8'h00}, /* 0xc287 */
            {8'h00}, /* 0xc286 */
            {8'h00}, /* 0xc285 */
            {8'h00}, /* 0xc284 */
            {8'h00}, /* 0xc283 */
            {8'h00}, /* 0xc282 */
            {8'h00}, /* 0xc281 */
            {8'h00}, /* 0xc280 */
            {8'h00}, /* 0xc27f */
            {8'h00}, /* 0xc27e */
            {8'h00}, /* 0xc27d */
            {8'h00}, /* 0xc27c */
            {8'h00}, /* 0xc27b */
            {8'h00}, /* 0xc27a */
            {8'h00}, /* 0xc279 */
            {8'h00}, /* 0xc278 */
            {8'h00}, /* 0xc277 */
            {8'h00}, /* 0xc276 */
            {8'h00}, /* 0xc275 */
            {8'h00}, /* 0xc274 */
            {8'h00}, /* 0xc273 */
            {8'h00}, /* 0xc272 */
            {8'h00}, /* 0xc271 */
            {8'h00}, /* 0xc270 */
            {8'h00}, /* 0xc26f */
            {8'h00}, /* 0xc26e */
            {8'h00}, /* 0xc26d */
            {8'h00}, /* 0xc26c */
            {8'h00}, /* 0xc26b */
            {8'h00}, /* 0xc26a */
            {8'h00}, /* 0xc269 */
            {8'h00}, /* 0xc268 */
            {8'h00}, /* 0xc267 */
            {8'h00}, /* 0xc266 */
            {8'h00}, /* 0xc265 */
            {8'h00}, /* 0xc264 */
            {8'h00}, /* 0xc263 */
            {8'h00}, /* 0xc262 */
            {8'h00}, /* 0xc261 */
            {8'h00}, /* 0xc260 */
            {8'h00}, /* 0xc25f */
            {8'h00}, /* 0xc25e */
            {8'h00}, /* 0xc25d */
            {8'h00}, /* 0xc25c */
            {8'h00}, /* 0xc25b */
            {8'h00}, /* 0xc25a */
            {8'h00}, /* 0xc259 */
            {8'h00}, /* 0xc258 */
            {8'h00}, /* 0xc257 */
            {8'h00}, /* 0xc256 */
            {8'h00}, /* 0xc255 */
            {8'h00}, /* 0xc254 */
            {8'h00}, /* 0xc253 */
            {8'h00}, /* 0xc252 */
            {8'h00}, /* 0xc251 */
            {8'h00}, /* 0xc250 */
            {8'h00}, /* 0xc24f */
            {8'h00}, /* 0xc24e */
            {8'h00}, /* 0xc24d */
            {8'h00}, /* 0xc24c */
            {8'h00}, /* 0xc24b */
            {8'h00}, /* 0xc24a */
            {8'h00}, /* 0xc249 */
            {8'h00}, /* 0xc248 */
            {8'h00}, /* 0xc247 */
            {8'h00}, /* 0xc246 */
            {8'h00}, /* 0xc245 */
            {8'h00}, /* 0xc244 */
            {8'h00}, /* 0xc243 */
            {8'h00}, /* 0xc242 */
            {8'h00}, /* 0xc241 */
            {8'h00}, /* 0xc240 */
            {8'h00}, /* 0xc23f */
            {8'h00}, /* 0xc23e */
            {8'h00}, /* 0xc23d */
            {8'h00}, /* 0xc23c */
            {8'h00}, /* 0xc23b */
            {8'h00}, /* 0xc23a */
            {8'h00}, /* 0xc239 */
            {8'h00}, /* 0xc238 */
            {8'h00}, /* 0xc237 */
            {8'h00}, /* 0xc236 */
            {8'h00}, /* 0xc235 */
            {8'h00}, /* 0xc234 */
            {8'h00}, /* 0xc233 */
            {8'h00}, /* 0xc232 */
            {8'h00}, /* 0xc231 */
            {8'h00}, /* 0xc230 */
            {8'h00}, /* 0xc22f */
            {8'h00}, /* 0xc22e */
            {8'h00}, /* 0xc22d */
            {8'h00}, /* 0xc22c */
            {8'h00}, /* 0xc22b */
            {8'h00}, /* 0xc22a */
            {8'h00}, /* 0xc229 */
            {8'h00}, /* 0xc228 */
            {8'h00}, /* 0xc227 */
            {8'h00}, /* 0xc226 */
            {8'h00}, /* 0xc225 */
            {8'h00}, /* 0xc224 */
            {8'h00}, /* 0xc223 */
            {8'h00}, /* 0xc222 */
            {8'h00}, /* 0xc221 */
            {8'h00}, /* 0xc220 */
            {8'h00}, /* 0xc21f */
            {8'h00}, /* 0xc21e */
            {8'h00}, /* 0xc21d */
            {8'h00}, /* 0xc21c */
            {8'h00}, /* 0xc21b */
            {8'h00}, /* 0xc21a */
            {8'h00}, /* 0xc219 */
            {8'h00}, /* 0xc218 */
            {8'h00}, /* 0xc217 */
            {8'h00}, /* 0xc216 */
            {8'h00}, /* 0xc215 */
            {8'h00}, /* 0xc214 */
            {8'h00}, /* 0xc213 */
            {8'h00}, /* 0xc212 */
            {8'h00}, /* 0xc211 */
            {8'h00}, /* 0xc210 */
            {8'h00}, /* 0xc20f */
            {8'h00}, /* 0xc20e */
            {8'h00}, /* 0xc20d */
            {8'h00}, /* 0xc20c */
            {8'h00}, /* 0xc20b */
            {8'h00}, /* 0xc20a */
            {8'h00}, /* 0xc209 */
            {8'h00}, /* 0xc208 */
            {8'h00}, /* 0xc207 */
            {8'h00}, /* 0xc206 */
            {8'h00}, /* 0xc205 */
            {8'h00}, /* 0xc204 */
            {8'h00}, /* 0xc203 */
            {8'h00}, /* 0xc202 */
            {8'h00}, /* 0xc201 */
            {8'h00}, /* 0xc200 */
            {8'h00}, /* 0xc1ff */
            {8'h00}, /* 0xc1fe */
            {8'h00}, /* 0xc1fd */
            {8'h00}, /* 0xc1fc */
            {8'h00}, /* 0xc1fb */
            {8'h00}, /* 0xc1fa */
            {8'h00}, /* 0xc1f9 */
            {8'h00}, /* 0xc1f8 */
            {8'h00}, /* 0xc1f7 */
            {8'h00}, /* 0xc1f6 */
            {8'h00}, /* 0xc1f5 */
            {8'h00}, /* 0xc1f4 */
            {8'h00}, /* 0xc1f3 */
            {8'h00}, /* 0xc1f2 */
            {8'h00}, /* 0xc1f1 */
            {8'h00}, /* 0xc1f0 */
            {8'h00}, /* 0xc1ef */
            {8'h00}, /* 0xc1ee */
            {8'h00}, /* 0xc1ed */
            {8'h00}, /* 0xc1ec */
            {8'h00}, /* 0xc1eb */
            {8'h00}, /* 0xc1ea */
            {8'h00}, /* 0xc1e9 */
            {8'h00}, /* 0xc1e8 */
            {8'h00}, /* 0xc1e7 */
            {8'h00}, /* 0xc1e6 */
            {8'h00}, /* 0xc1e5 */
            {8'h00}, /* 0xc1e4 */
            {8'h00}, /* 0xc1e3 */
            {8'h00}, /* 0xc1e2 */
            {8'h00}, /* 0xc1e1 */
            {8'h00}, /* 0xc1e0 */
            {8'h00}, /* 0xc1df */
            {8'h00}, /* 0xc1de */
            {8'h00}, /* 0xc1dd */
            {8'h00}, /* 0xc1dc */
            {8'h00}, /* 0xc1db */
            {8'h00}, /* 0xc1da */
            {8'h00}, /* 0xc1d9 */
            {8'h00}, /* 0xc1d8 */
            {8'h00}, /* 0xc1d7 */
            {8'h00}, /* 0xc1d6 */
            {8'h00}, /* 0xc1d5 */
            {8'h00}, /* 0xc1d4 */
            {8'h00}, /* 0xc1d3 */
            {8'h00}, /* 0xc1d2 */
            {8'h00}, /* 0xc1d1 */
            {8'h00}, /* 0xc1d0 */
            {8'h00}, /* 0xc1cf */
            {8'h00}, /* 0xc1ce */
            {8'h00}, /* 0xc1cd */
            {8'h00}, /* 0xc1cc */
            {8'h00}, /* 0xc1cb */
            {8'h00}, /* 0xc1ca */
            {8'h00}, /* 0xc1c9 */
            {8'h00}, /* 0xc1c8 */
            {8'h00}, /* 0xc1c7 */
            {8'h00}, /* 0xc1c6 */
            {8'h00}, /* 0xc1c5 */
            {8'h00}, /* 0xc1c4 */
            {8'h00}, /* 0xc1c3 */
            {8'h00}, /* 0xc1c2 */
            {8'h00}, /* 0xc1c1 */
            {8'h00}, /* 0xc1c0 */
            {8'h00}, /* 0xc1bf */
            {8'h00}, /* 0xc1be */
            {8'h00}, /* 0xc1bd */
            {8'h00}, /* 0xc1bc */
            {8'h00}, /* 0xc1bb */
            {8'h00}, /* 0xc1ba */
            {8'h00}, /* 0xc1b9 */
            {8'h00}, /* 0xc1b8 */
            {8'h00}, /* 0xc1b7 */
            {8'h00}, /* 0xc1b6 */
            {8'h00}, /* 0xc1b5 */
            {8'h00}, /* 0xc1b4 */
            {8'h00}, /* 0xc1b3 */
            {8'h00}, /* 0xc1b2 */
            {8'h00}, /* 0xc1b1 */
            {8'h00}, /* 0xc1b0 */
            {8'h00}, /* 0xc1af */
            {8'h00}, /* 0xc1ae */
            {8'h00}, /* 0xc1ad */
            {8'h00}, /* 0xc1ac */
            {8'h00}, /* 0xc1ab */
            {8'h00}, /* 0xc1aa */
            {8'h00}, /* 0xc1a9 */
            {8'h00}, /* 0xc1a8 */
            {8'h00}, /* 0xc1a7 */
            {8'h00}, /* 0xc1a6 */
            {8'h00}, /* 0xc1a5 */
            {8'h00}, /* 0xc1a4 */
            {8'h00}, /* 0xc1a3 */
            {8'h00}, /* 0xc1a2 */
            {8'h00}, /* 0xc1a1 */
            {8'h00}, /* 0xc1a0 */
            {8'h00}, /* 0xc19f */
            {8'h00}, /* 0xc19e */
            {8'h00}, /* 0xc19d */
            {8'h00}, /* 0xc19c */
            {8'h00}, /* 0xc19b */
            {8'h00}, /* 0xc19a */
            {8'h00}, /* 0xc199 */
            {8'h00}, /* 0xc198 */
            {8'h00}, /* 0xc197 */
            {8'h00}, /* 0xc196 */
            {8'h00}, /* 0xc195 */
            {8'h00}, /* 0xc194 */
            {8'h00}, /* 0xc193 */
            {8'h00}, /* 0xc192 */
            {8'h00}, /* 0xc191 */
            {8'h00}, /* 0xc190 */
            {8'h00}, /* 0xc18f */
            {8'h00}, /* 0xc18e */
            {8'h00}, /* 0xc18d */
            {8'h00}, /* 0xc18c */
            {8'h00}, /* 0xc18b */
            {8'h00}, /* 0xc18a */
            {8'h00}, /* 0xc189 */
            {8'h00}, /* 0xc188 */
            {8'h00}, /* 0xc187 */
            {8'h00}, /* 0xc186 */
            {8'h00}, /* 0xc185 */
            {8'h00}, /* 0xc184 */
            {8'h00}, /* 0xc183 */
            {8'h00}, /* 0xc182 */
            {8'h00}, /* 0xc181 */
            {8'h00}, /* 0xc180 */
            {8'h00}, /* 0xc17f */
            {8'h00}, /* 0xc17e */
            {8'h00}, /* 0xc17d */
            {8'h00}, /* 0xc17c */
            {8'h00}, /* 0xc17b */
            {8'h00}, /* 0xc17a */
            {8'h00}, /* 0xc179 */
            {8'h00}, /* 0xc178 */
            {8'h00}, /* 0xc177 */
            {8'h00}, /* 0xc176 */
            {8'h00}, /* 0xc175 */
            {8'h00}, /* 0xc174 */
            {8'h00}, /* 0xc173 */
            {8'h00}, /* 0xc172 */
            {8'h00}, /* 0xc171 */
            {8'h00}, /* 0xc170 */
            {8'h00}, /* 0xc16f */
            {8'h00}, /* 0xc16e */
            {8'h00}, /* 0xc16d */
            {8'h00}, /* 0xc16c */
            {8'h00}, /* 0xc16b */
            {8'h00}, /* 0xc16a */
            {8'h00}, /* 0xc169 */
            {8'h00}, /* 0xc168 */
            {8'h00}, /* 0xc167 */
            {8'h00}, /* 0xc166 */
            {8'h00}, /* 0xc165 */
            {8'h00}, /* 0xc164 */
            {8'h00}, /* 0xc163 */
            {8'h00}, /* 0xc162 */
            {8'h00}, /* 0xc161 */
            {8'h00}, /* 0xc160 */
            {8'h00}, /* 0xc15f */
            {8'h00}, /* 0xc15e */
            {8'h00}, /* 0xc15d */
            {8'h00}, /* 0xc15c */
            {8'h00}, /* 0xc15b */
            {8'h00}, /* 0xc15a */
            {8'h00}, /* 0xc159 */
            {8'h00}, /* 0xc158 */
            {8'h00}, /* 0xc157 */
            {8'h00}, /* 0xc156 */
            {8'h00}, /* 0xc155 */
            {8'h00}, /* 0xc154 */
            {8'h00}, /* 0xc153 */
            {8'h00}, /* 0xc152 */
            {8'h00}, /* 0xc151 */
            {8'h00}, /* 0xc150 */
            {8'h00}, /* 0xc14f */
            {8'h00}, /* 0xc14e */
            {8'h00}, /* 0xc14d */
            {8'h00}, /* 0xc14c */
            {8'h00}, /* 0xc14b */
            {8'h00}, /* 0xc14a */
            {8'h00}, /* 0xc149 */
            {8'h00}, /* 0xc148 */
            {8'h00}, /* 0xc147 */
            {8'h00}, /* 0xc146 */
            {8'h00}, /* 0xc145 */
            {8'h00}, /* 0xc144 */
            {8'h00}, /* 0xc143 */
            {8'h00}, /* 0xc142 */
            {8'h00}, /* 0xc141 */
            {8'h00}, /* 0xc140 */
            {8'h00}, /* 0xc13f */
            {8'h00}, /* 0xc13e */
            {8'h00}, /* 0xc13d */
            {8'h00}, /* 0xc13c */
            {8'h00}, /* 0xc13b */
            {8'h00}, /* 0xc13a */
            {8'h00}, /* 0xc139 */
            {8'h00}, /* 0xc138 */
            {8'h00}, /* 0xc137 */
            {8'h00}, /* 0xc136 */
            {8'h00}, /* 0xc135 */
            {8'h00}, /* 0xc134 */
            {8'h00}, /* 0xc133 */
            {8'h00}, /* 0xc132 */
            {8'h00}, /* 0xc131 */
            {8'h00}, /* 0xc130 */
            {8'h00}, /* 0xc12f */
            {8'h00}, /* 0xc12e */
            {8'h00}, /* 0xc12d */
            {8'h00}, /* 0xc12c */
            {8'h00}, /* 0xc12b */
            {8'h00}, /* 0xc12a */
            {8'h00}, /* 0xc129 */
            {8'h00}, /* 0xc128 */
            {8'h00}, /* 0xc127 */
            {8'h00}, /* 0xc126 */
            {8'h00}, /* 0xc125 */
            {8'h00}, /* 0xc124 */
            {8'h00}, /* 0xc123 */
            {8'h00}, /* 0xc122 */
            {8'h00}, /* 0xc121 */
            {8'h00}, /* 0xc120 */
            {8'h00}, /* 0xc11f */
            {8'h00}, /* 0xc11e */
            {8'h00}, /* 0xc11d */
            {8'h00}, /* 0xc11c */
            {8'h00}, /* 0xc11b */
            {8'h00}, /* 0xc11a */
            {8'h00}, /* 0xc119 */
            {8'h00}, /* 0xc118 */
            {8'h00}, /* 0xc117 */
            {8'h00}, /* 0xc116 */
            {8'h00}, /* 0xc115 */
            {8'h00}, /* 0xc114 */
            {8'h00}, /* 0xc113 */
            {8'h00}, /* 0xc112 */
            {8'h00}, /* 0xc111 */
            {8'h00}, /* 0xc110 */
            {8'h00}, /* 0xc10f */
            {8'h00}, /* 0xc10e */
            {8'h00}, /* 0xc10d */
            {8'h00}, /* 0xc10c */
            {8'h00}, /* 0xc10b */
            {8'h00}, /* 0xc10a */
            {8'h00}, /* 0xc109 */
            {8'h00}, /* 0xc108 */
            {8'h00}, /* 0xc107 */
            {8'h00}, /* 0xc106 */
            {8'h00}, /* 0xc105 */
            {8'h00}, /* 0xc104 */
            {8'h00}, /* 0xc103 */
            {8'h00}, /* 0xc102 */
            {8'h00}, /* 0xc101 */
            {8'h00}, /* 0xc100 */
            {8'h00}, /* 0xc0ff */
            {8'h00}, /* 0xc0fe */
            {8'h00}, /* 0xc0fd */
            {8'h00}, /* 0xc0fc */
            {8'h00}, /* 0xc0fb */
            {8'h00}, /* 0xc0fa */
            {8'h00}, /* 0xc0f9 */
            {8'h00}, /* 0xc0f8 */
            {8'h00}, /* 0xc0f7 */
            {8'h00}, /* 0xc0f6 */
            {8'h00}, /* 0xc0f5 */
            {8'h00}, /* 0xc0f4 */
            {8'h00}, /* 0xc0f3 */
            {8'h00}, /* 0xc0f2 */
            {8'h00}, /* 0xc0f1 */
            {8'h00}, /* 0xc0f0 */
            {8'h00}, /* 0xc0ef */
            {8'h00}, /* 0xc0ee */
            {8'h00}, /* 0xc0ed */
            {8'h00}, /* 0xc0ec */
            {8'h00}, /* 0xc0eb */
            {8'h00}, /* 0xc0ea */
            {8'h00}, /* 0xc0e9 */
            {8'h00}, /* 0xc0e8 */
            {8'h00}, /* 0xc0e7 */
            {8'h00}, /* 0xc0e6 */
            {8'h00}, /* 0xc0e5 */
            {8'h00}, /* 0xc0e4 */
            {8'h00}, /* 0xc0e3 */
            {8'h00}, /* 0xc0e2 */
            {8'h00}, /* 0xc0e1 */
            {8'h00}, /* 0xc0e0 */
            {8'h00}, /* 0xc0df */
            {8'h00}, /* 0xc0de */
            {8'h00}, /* 0xc0dd */
            {8'h00}, /* 0xc0dc */
            {8'h00}, /* 0xc0db */
            {8'h00}, /* 0xc0da */
            {8'h00}, /* 0xc0d9 */
            {8'h00}, /* 0xc0d8 */
            {8'h00}, /* 0xc0d7 */
            {8'h00}, /* 0xc0d6 */
            {8'h00}, /* 0xc0d5 */
            {8'h00}, /* 0xc0d4 */
            {8'h00}, /* 0xc0d3 */
            {8'h00}, /* 0xc0d2 */
            {8'h00}, /* 0xc0d1 */
            {8'h00}, /* 0xc0d0 */
            {8'h00}, /* 0xc0cf */
            {8'h00}, /* 0xc0ce */
            {8'h00}, /* 0xc0cd */
            {8'h00}, /* 0xc0cc */
            {8'h00}, /* 0xc0cb */
            {8'h00}, /* 0xc0ca */
            {8'h00}, /* 0xc0c9 */
            {8'h00}, /* 0xc0c8 */
            {8'h00}, /* 0xc0c7 */
            {8'h00}, /* 0xc0c6 */
            {8'h00}, /* 0xc0c5 */
            {8'h00}, /* 0xc0c4 */
            {8'h00}, /* 0xc0c3 */
            {8'h00}, /* 0xc0c2 */
            {8'h00}, /* 0xc0c1 */
            {8'h00}, /* 0xc0c0 */
            {8'h00}, /* 0xc0bf */
            {8'h00}, /* 0xc0be */
            {8'h00}, /* 0xc0bd */
            {8'h00}, /* 0xc0bc */
            {8'h00}, /* 0xc0bb */
            {8'h00}, /* 0xc0ba */
            {8'h00}, /* 0xc0b9 */
            {8'h00}, /* 0xc0b8 */
            {8'h00}, /* 0xc0b7 */
            {8'h00}, /* 0xc0b6 */
            {8'h00}, /* 0xc0b5 */
            {8'h00}, /* 0xc0b4 */
            {8'h00}, /* 0xc0b3 */
            {8'h00}, /* 0xc0b2 */
            {8'h00}, /* 0xc0b1 */
            {8'h00}, /* 0xc0b0 */
            {8'h00}, /* 0xc0af */
            {8'h00}, /* 0xc0ae */
            {8'h00}, /* 0xc0ad */
            {8'h00}, /* 0xc0ac */
            {8'h00}, /* 0xc0ab */
            {8'h00}, /* 0xc0aa */
            {8'h00}, /* 0xc0a9 */
            {8'h00}, /* 0xc0a8 */
            {8'h00}, /* 0xc0a7 */
            {8'h00}, /* 0xc0a6 */
            {8'h00}, /* 0xc0a5 */
            {8'h00}, /* 0xc0a4 */
            {8'h00}, /* 0xc0a3 */
            {8'h00}, /* 0xc0a2 */
            {8'h00}, /* 0xc0a1 */
            {8'h00}, /* 0xc0a0 */
            {8'h00}, /* 0xc09f */
            {8'h00}, /* 0xc09e */
            {8'h00}, /* 0xc09d */
            {8'h00}, /* 0xc09c */
            {8'h00}, /* 0xc09b */
            {8'h00}, /* 0xc09a */
            {8'h00}, /* 0xc099 */
            {8'h00}, /* 0xc098 */
            {8'h00}, /* 0xc097 */
            {8'h00}, /* 0xc096 */
            {8'h00}, /* 0xc095 */
            {8'h00}, /* 0xc094 */
            {8'h00}, /* 0xc093 */
            {8'h00}, /* 0xc092 */
            {8'h00}, /* 0xc091 */
            {8'h00}, /* 0xc090 */
            {8'h00}, /* 0xc08f */
            {8'h00}, /* 0xc08e */
            {8'h00}, /* 0xc08d */
            {8'h00}, /* 0xc08c */
            {8'h00}, /* 0xc08b */
            {8'h00}, /* 0xc08a */
            {8'h00}, /* 0xc089 */
            {8'h00}, /* 0xc088 */
            {8'h00}, /* 0xc087 */
            {8'h00}, /* 0xc086 */
            {8'h00}, /* 0xc085 */
            {8'h00}, /* 0xc084 */
            {8'h00}, /* 0xc083 */
            {8'h00}, /* 0xc082 */
            {8'h00}, /* 0xc081 */
            {8'h00}, /* 0xc080 */
            {8'h00}, /* 0xc07f */
            {8'h00}, /* 0xc07e */
            {8'h00}, /* 0xc07d */
            {8'h00}, /* 0xc07c */
            {8'h00}, /* 0xc07b */
            {8'h00}, /* 0xc07a */
            {8'h00}, /* 0xc079 */
            {8'h00}, /* 0xc078 */
            {8'h00}, /* 0xc077 */
            {8'h00}, /* 0xc076 */
            {8'h00}, /* 0xc075 */
            {8'h00}, /* 0xc074 */
            {8'h00}, /* 0xc073 */
            {8'h00}, /* 0xc072 */
            {8'h00}, /* 0xc071 */
            {8'h00}, /* 0xc070 */
            {8'h00}, /* 0xc06f */
            {8'h00}, /* 0xc06e */
            {8'h00}, /* 0xc06d */
            {8'h00}, /* 0xc06c */
            {8'h00}, /* 0xc06b */
            {8'h00}, /* 0xc06a */
            {8'h00}, /* 0xc069 */
            {8'h00}, /* 0xc068 */
            {8'h00}, /* 0xc067 */
            {8'h00}, /* 0xc066 */
            {8'h00}, /* 0xc065 */
            {8'h00}, /* 0xc064 */
            {8'h00}, /* 0xc063 */
            {8'h00}, /* 0xc062 */
            {8'h00}, /* 0xc061 */
            {8'h00}, /* 0xc060 */
            {8'h00}, /* 0xc05f */
            {8'h00}, /* 0xc05e */
            {8'h00}, /* 0xc05d */
            {8'h00}, /* 0xc05c */
            {8'h00}, /* 0xc05b */
            {8'h00}, /* 0xc05a */
            {8'h00}, /* 0xc059 */
            {8'h00}, /* 0xc058 */
            {8'h00}, /* 0xc057 */
            {8'h00}, /* 0xc056 */
            {8'h00}, /* 0xc055 */
            {8'h00}, /* 0xc054 */
            {8'h00}, /* 0xc053 */
            {8'h00}, /* 0xc052 */
            {8'h00}, /* 0xc051 */
            {8'h00}, /* 0xc050 */
            {8'h00}, /* 0xc04f */
            {8'h00}, /* 0xc04e */
            {8'h00}, /* 0xc04d */
            {8'h00}, /* 0xc04c */
            {8'h00}, /* 0xc04b */
            {8'h00}, /* 0xc04a */
            {8'h00}, /* 0xc049 */
            {8'h00}, /* 0xc048 */
            {8'h00}, /* 0xc047 */
            {8'h00}, /* 0xc046 */
            {8'h00}, /* 0xc045 */
            {8'h00}, /* 0xc044 */
            {8'h00}, /* 0xc043 */
            {8'h00}, /* 0xc042 */
            {8'h00}, /* 0xc041 */
            {8'h00}, /* 0xc040 */
            {8'h00}, /* 0xc03f */
            {8'h00}, /* 0xc03e */
            {8'h00}, /* 0xc03d */
            {8'h00}, /* 0xc03c */
            {8'h00}, /* 0xc03b */
            {8'h00}, /* 0xc03a */
            {8'h00}, /* 0xc039 */
            {8'h00}, /* 0xc038 */
            {8'h00}, /* 0xc037 */
            {8'h00}, /* 0xc036 */
            {8'h00}, /* 0xc035 */
            {8'h00}, /* 0xc034 */
            {8'h00}, /* 0xc033 */
            {8'h00}, /* 0xc032 */
            {8'h00}, /* 0xc031 */
            {8'h00}, /* 0xc030 */
            {8'h00}, /* 0xc02f */
            {8'h00}, /* 0xc02e */
            {8'h00}, /* 0xc02d */
            {8'h00}, /* 0xc02c */
            {8'h00}, /* 0xc02b */
            {8'h00}, /* 0xc02a */
            {8'h00}, /* 0xc029 */
            {8'h00}, /* 0xc028 */
            {8'h00}, /* 0xc027 */
            {8'h00}, /* 0xc026 */
            {8'h00}, /* 0xc025 */
            {8'h00}, /* 0xc024 */
            {8'h00}, /* 0xc023 */
            {8'h00}, /* 0xc022 */
            {8'h00}, /* 0xc021 */
            {8'h00}, /* 0xc020 */
            {8'h00}, /* 0xc01f */
            {8'h00}, /* 0xc01e */
            {8'h00}, /* 0xc01d */
            {8'h00}, /* 0xc01c */
            {8'h00}, /* 0xc01b */
            {8'h00}, /* 0xc01a */
            {8'h00}, /* 0xc019 */
            {8'h00}, /* 0xc018 */
            {8'h00}, /* 0xc017 */
            {8'h00}, /* 0xc016 */
            {8'h00}, /* 0xc015 */
            {8'h00}, /* 0xc014 */
            {8'h00}, /* 0xc013 */
            {8'h00}, /* 0xc012 */
            {8'h00}, /* 0xc011 */
            {8'h00}, /* 0xc010 */
            {8'h00}, /* 0xc00f */
            {8'h00}, /* 0xc00e */
            {8'h00}, /* 0xc00d */
            {8'h00}, /* 0xc00c */
            {8'h00}, /* 0xc00b */
            {8'h00}, /* 0xc00a */
            {8'h00}, /* 0xc009 */
            {8'h00}, /* 0xc008 */
            {8'h00}, /* 0xc007 */
            {8'h00}, /* 0xc006 */
            {8'h00}, /* 0xc005 */
            {8'h00}, /* 0xc004 */
            {8'h00}, /* 0xc003 */
            {8'h00}, /* 0xc002 */
            {8'h00}, /* 0xc001 */
            {8'h00}, /* 0xc000 */
            {8'h00}, /* 0xbfff */
            {8'h00}, /* 0xbffe */
            {8'h00}, /* 0xbffd */
            {8'h00}, /* 0xbffc */
            {8'h00}, /* 0xbffb */
            {8'h00}, /* 0xbffa */
            {8'h00}, /* 0xbff9 */
            {8'h00}, /* 0xbff8 */
            {8'h00}, /* 0xbff7 */
            {8'h00}, /* 0xbff6 */
            {8'h00}, /* 0xbff5 */
            {8'h00}, /* 0xbff4 */
            {8'h00}, /* 0xbff3 */
            {8'h00}, /* 0xbff2 */
            {8'h00}, /* 0xbff1 */
            {8'h00}, /* 0xbff0 */
            {8'h00}, /* 0xbfef */
            {8'h00}, /* 0xbfee */
            {8'h00}, /* 0xbfed */
            {8'h00}, /* 0xbfec */
            {8'h00}, /* 0xbfeb */
            {8'h00}, /* 0xbfea */
            {8'h00}, /* 0xbfe9 */
            {8'h00}, /* 0xbfe8 */
            {8'h00}, /* 0xbfe7 */
            {8'h00}, /* 0xbfe6 */
            {8'h00}, /* 0xbfe5 */
            {8'h00}, /* 0xbfe4 */
            {8'h00}, /* 0xbfe3 */
            {8'h00}, /* 0xbfe2 */
            {8'h00}, /* 0xbfe1 */
            {8'h00}, /* 0xbfe0 */
            {8'h00}, /* 0xbfdf */
            {8'h00}, /* 0xbfde */
            {8'h00}, /* 0xbfdd */
            {8'h00}, /* 0xbfdc */
            {8'h00}, /* 0xbfdb */
            {8'h00}, /* 0xbfda */
            {8'h00}, /* 0xbfd9 */
            {8'h00}, /* 0xbfd8 */
            {8'h00}, /* 0xbfd7 */
            {8'h00}, /* 0xbfd6 */
            {8'h00}, /* 0xbfd5 */
            {8'h00}, /* 0xbfd4 */
            {8'h00}, /* 0xbfd3 */
            {8'h00}, /* 0xbfd2 */
            {8'h00}, /* 0xbfd1 */
            {8'h00}, /* 0xbfd0 */
            {8'h00}, /* 0xbfcf */
            {8'h00}, /* 0xbfce */
            {8'h00}, /* 0xbfcd */
            {8'h00}, /* 0xbfcc */
            {8'h00}, /* 0xbfcb */
            {8'h00}, /* 0xbfca */
            {8'h00}, /* 0xbfc9 */
            {8'h00}, /* 0xbfc8 */
            {8'h00}, /* 0xbfc7 */
            {8'h00}, /* 0xbfc6 */
            {8'h00}, /* 0xbfc5 */
            {8'h00}, /* 0xbfc4 */
            {8'h00}, /* 0xbfc3 */
            {8'h00}, /* 0xbfc2 */
            {8'h00}, /* 0xbfc1 */
            {8'h00}, /* 0xbfc0 */
            {8'h00}, /* 0xbfbf */
            {8'h00}, /* 0xbfbe */
            {8'h00}, /* 0xbfbd */
            {8'h00}, /* 0xbfbc */
            {8'h00}, /* 0xbfbb */
            {8'h00}, /* 0xbfba */
            {8'h00}, /* 0xbfb9 */
            {8'h00}, /* 0xbfb8 */
            {8'h00}, /* 0xbfb7 */
            {8'h00}, /* 0xbfb6 */
            {8'h00}, /* 0xbfb5 */
            {8'h00}, /* 0xbfb4 */
            {8'h00}, /* 0xbfb3 */
            {8'h00}, /* 0xbfb2 */
            {8'h00}, /* 0xbfb1 */
            {8'h00}, /* 0xbfb0 */
            {8'h00}, /* 0xbfaf */
            {8'h00}, /* 0xbfae */
            {8'h00}, /* 0xbfad */
            {8'h00}, /* 0xbfac */
            {8'h00}, /* 0xbfab */
            {8'h00}, /* 0xbfaa */
            {8'h00}, /* 0xbfa9 */
            {8'h00}, /* 0xbfa8 */
            {8'h00}, /* 0xbfa7 */
            {8'h00}, /* 0xbfa6 */
            {8'h00}, /* 0xbfa5 */
            {8'h00}, /* 0xbfa4 */
            {8'h00}, /* 0xbfa3 */
            {8'h00}, /* 0xbfa2 */
            {8'h00}, /* 0xbfa1 */
            {8'h00}, /* 0xbfa0 */
            {8'h00}, /* 0xbf9f */
            {8'h00}, /* 0xbf9e */
            {8'h00}, /* 0xbf9d */
            {8'h00}, /* 0xbf9c */
            {8'h00}, /* 0xbf9b */
            {8'h00}, /* 0xbf9a */
            {8'h00}, /* 0xbf99 */
            {8'h00}, /* 0xbf98 */
            {8'h00}, /* 0xbf97 */
            {8'h00}, /* 0xbf96 */
            {8'h00}, /* 0xbf95 */
            {8'h00}, /* 0xbf94 */
            {8'h00}, /* 0xbf93 */
            {8'h00}, /* 0xbf92 */
            {8'h00}, /* 0xbf91 */
            {8'h00}, /* 0xbf90 */
            {8'h00}, /* 0xbf8f */
            {8'h00}, /* 0xbf8e */
            {8'h00}, /* 0xbf8d */
            {8'h00}, /* 0xbf8c */
            {8'h00}, /* 0xbf8b */
            {8'h00}, /* 0xbf8a */
            {8'h00}, /* 0xbf89 */
            {8'h00}, /* 0xbf88 */
            {8'h00}, /* 0xbf87 */
            {8'h00}, /* 0xbf86 */
            {8'h00}, /* 0xbf85 */
            {8'h00}, /* 0xbf84 */
            {8'h00}, /* 0xbf83 */
            {8'h00}, /* 0xbf82 */
            {8'h00}, /* 0xbf81 */
            {8'h00}, /* 0xbf80 */
            {8'h00}, /* 0xbf7f */
            {8'h00}, /* 0xbf7e */
            {8'h00}, /* 0xbf7d */
            {8'h00}, /* 0xbf7c */
            {8'h00}, /* 0xbf7b */
            {8'h00}, /* 0xbf7a */
            {8'h00}, /* 0xbf79 */
            {8'h00}, /* 0xbf78 */
            {8'h00}, /* 0xbf77 */
            {8'h00}, /* 0xbf76 */
            {8'h00}, /* 0xbf75 */
            {8'h00}, /* 0xbf74 */
            {8'h00}, /* 0xbf73 */
            {8'h00}, /* 0xbf72 */
            {8'h00}, /* 0xbf71 */
            {8'h00}, /* 0xbf70 */
            {8'h00}, /* 0xbf6f */
            {8'h00}, /* 0xbf6e */
            {8'h00}, /* 0xbf6d */
            {8'h00}, /* 0xbf6c */
            {8'h00}, /* 0xbf6b */
            {8'h00}, /* 0xbf6a */
            {8'h00}, /* 0xbf69 */
            {8'h00}, /* 0xbf68 */
            {8'h00}, /* 0xbf67 */
            {8'h00}, /* 0xbf66 */
            {8'h00}, /* 0xbf65 */
            {8'h00}, /* 0xbf64 */
            {8'h00}, /* 0xbf63 */
            {8'h00}, /* 0xbf62 */
            {8'h00}, /* 0xbf61 */
            {8'h00}, /* 0xbf60 */
            {8'h00}, /* 0xbf5f */
            {8'h00}, /* 0xbf5e */
            {8'h00}, /* 0xbf5d */
            {8'h00}, /* 0xbf5c */
            {8'h00}, /* 0xbf5b */
            {8'h00}, /* 0xbf5a */
            {8'h00}, /* 0xbf59 */
            {8'h00}, /* 0xbf58 */
            {8'h00}, /* 0xbf57 */
            {8'h00}, /* 0xbf56 */
            {8'h00}, /* 0xbf55 */
            {8'h00}, /* 0xbf54 */
            {8'h00}, /* 0xbf53 */
            {8'h00}, /* 0xbf52 */
            {8'h00}, /* 0xbf51 */
            {8'h00}, /* 0xbf50 */
            {8'h00}, /* 0xbf4f */
            {8'h00}, /* 0xbf4e */
            {8'h00}, /* 0xbf4d */
            {8'h00}, /* 0xbf4c */
            {8'h00}, /* 0xbf4b */
            {8'h00}, /* 0xbf4a */
            {8'h00}, /* 0xbf49 */
            {8'h00}, /* 0xbf48 */
            {8'h00}, /* 0xbf47 */
            {8'h00}, /* 0xbf46 */
            {8'h00}, /* 0xbf45 */
            {8'h00}, /* 0xbf44 */
            {8'h00}, /* 0xbf43 */
            {8'h00}, /* 0xbf42 */
            {8'h00}, /* 0xbf41 */
            {8'h00}, /* 0xbf40 */
            {8'h00}, /* 0xbf3f */
            {8'h00}, /* 0xbf3e */
            {8'h00}, /* 0xbf3d */
            {8'h00}, /* 0xbf3c */
            {8'h00}, /* 0xbf3b */
            {8'h00}, /* 0xbf3a */
            {8'h00}, /* 0xbf39 */
            {8'h00}, /* 0xbf38 */
            {8'h00}, /* 0xbf37 */
            {8'h00}, /* 0xbf36 */
            {8'h00}, /* 0xbf35 */
            {8'h00}, /* 0xbf34 */
            {8'h00}, /* 0xbf33 */
            {8'h00}, /* 0xbf32 */
            {8'h00}, /* 0xbf31 */
            {8'h00}, /* 0xbf30 */
            {8'h00}, /* 0xbf2f */
            {8'h00}, /* 0xbf2e */
            {8'h00}, /* 0xbf2d */
            {8'h00}, /* 0xbf2c */
            {8'h00}, /* 0xbf2b */
            {8'h00}, /* 0xbf2a */
            {8'h00}, /* 0xbf29 */
            {8'h00}, /* 0xbf28 */
            {8'h00}, /* 0xbf27 */
            {8'h00}, /* 0xbf26 */
            {8'h00}, /* 0xbf25 */
            {8'h00}, /* 0xbf24 */
            {8'h00}, /* 0xbf23 */
            {8'h00}, /* 0xbf22 */
            {8'h00}, /* 0xbf21 */
            {8'h00}, /* 0xbf20 */
            {8'h00}, /* 0xbf1f */
            {8'h00}, /* 0xbf1e */
            {8'h00}, /* 0xbf1d */
            {8'h00}, /* 0xbf1c */
            {8'h00}, /* 0xbf1b */
            {8'h00}, /* 0xbf1a */
            {8'h00}, /* 0xbf19 */
            {8'h00}, /* 0xbf18 */
            {8'h00}, /* 0xbf17 */
            {8'h00}, /* 0xbf16 */
            {8'h00}, /* 0xbf15 */
            {8'h00}, /* 0xbf14 */
            {8'h00}, /* 0xbf13 */
            {8'h00}, /* 0xbf12 */
            {8'h00}, /* 0xbf11 */
            {8'h00}, /* 0xbf10 */
            {8'h00}, /* 0xbf0f */
            {8'h00}, /* 0xbf0e */
            {8'h00}, /* 0xbf0d */
            {8'h00}, /* 0xbf0c */
            {8'h00}, /* 0xbf0b */
            {8'h00}, /* 0xbf0a */
            {8'h00}, /* 0xbf09 */
            {8'h00}, /* 0xbf08 */
            {8'h00}, /* 0xbf07 */
            {8'h00}, /* 0xbf06 */
            {8'h00}, /* 0xbf05 */
            {8'h00}, /* 0xbf04 */
            {8'h00}, /* 0xbf03 */
            {8'h00}, /* 0xbf02 */
            {8'h00}, /* 0xbf01 */
            {8'h00}, /* 0xbf00 */
            {8'h00}, /* 0xbeff */
            {8'h00}, /* 0xbefe */
            {8'h00}, /* 0xbefd */
            {8'h00}, /* 0xbefc */
            {8'h00}, /* 0xbefb */
            {8'h00}, /* 0xbefa */
            {8'h00}, /* 0xbef9 */
            {8'h00}, /* 0xbef8 */
            {8'h00}, /* 0xbef7 */
            {8'h00}, /* 0xbef6 */
            {8'h00}, /* 0xbef5 */
            {8'h00}, /* 0xbef4 */
            {8'h00}, /* 0xbef3 */
            {8'h00}, /* 0xbef2 */
            {8'h00}, /* 0xbef1 */
            {8'h00}, /* 0xbef0 */
            {8'h00}, /* 0xbeef */
            {8'h00}, /* 0xbeee */
            {8'h00}, /* 0xbeed */
            {8'h00}, /* 0xbeec */
            {8'h00}, /* 0xbeeb */
            {8'h00}, /* 0xbeea */
            {8'h00}, /* 0xbee9 */
            {8'h00}, /* 0xbee8 */
            {8'h00}, /* 0xbee7 */
            {8'h00}, /* 0xbee6 */
            {8'h00}, /* 0xbee5 */
            {8'h00}, /* 0xbee4 */
            {8'h00}, /* 0xbee3 */
            {8'h00}, /* 0xbee2 */
            {8'h00}, /* 0xbee1 */
            {8'h00}, /* 0xbee0 */
            {8'h00}, /* 0xbedf */
            {8'h00}, /* 0xbede */
            {8'h00}, /* 0xbedd */
            {8'h00}, /* 0xbedc */
            {8'h00}, /* 0xbedb */
            {8'h00}, /* 0xbeda */
            {8'h00}, /* 0xbed9 */
            {8'h00}, /* 0xbed8 */
            {8'h00}, /* 0xbed7 */
            {8'h00}, /* 0xbed6 */
            {8'h00}, /* 0xbed5 */
            {8'h00}, /* 0xbed4 */
            {8'h00}, /* 0xbed3 */
            {8'h00}, /* 0xbed2 */
            {8'h00}, /* 0xbed1 */
            {8'h00}, /* 0xbed0 */
            {8'h00}, /* 0xbecf */
            {8'h00}, /* 0xbece */
            {8'h00}, /* 0xbecd */
            {8'h00}, /* 0xbecc */
            {8'h00}, /* 0xbecb */
            {8'h00}, /* 0xbeca */
            {8'h00}, /* 0xbec9 */
            {8'h00}, /* 0xbec8 */
            {8'h00}, /* 0xbec7 */
            {8'h00}, /* 0xbec6 */
            {8'h00}, /* 0xbec5 */
            {8'h00}, /* 0xbec4 */
            {8'h00}, /* 0xbec3 */
            {8'h00}, /* 0xbec2 */
            {8'h00}, /* 0xbec1 */
            {8'h00}, /* 0xbec0 */
            {8'h00}, /* 0xbebf */
            {8'h00}, /* 0xbebe */
            {8'h00}, /* 0xbebd */
            {8'h00}, /* 0xbebc */
            {8'h00}, /* 0xbebb */
            {8'h00}, /* 0xbeba */
            {8'h00}, /* 0xbeb9 */
            {8'h00}, /* 0xbeb8 */
            {8'h00}, /* 0xbeb7 */
            {8'h00}, /* 0xbeb6 */
            {8'h00}, /* 0xbeb5 */
            {8'h00}, /* 0xbeb4 */
            {8'h00}, /* 0xbeb3 */
            {8'h00}, /* 0xbeb2 */
            {8'h00}, /* 0xbeb1 */
            {8'h00}, /* 0xbeb0 */
            {8'h00}, /* 0xbeaf */
            {8'h00}, /* 0xbeae */
            {8'h00}, /* 0xbead */
            {8'h00}, /* 0xbeac */
            {8'h00}, /* 0xbeab */
            {8'h00}, /* 0xbeaa */
            {8'h00}, /* 0xbea9 */
            {8'h00}, /* 0xbea8 */
            {8'h00}, /* 0xbea7 */
            {8'h00}, /* 0xbea6 */
            {8'h00}, /* 0xbea5 */
            {8'h00}, /* 0xbea4 */
            {8'h00}, /* 0xbea3 */
            {8'h00}, /* 0xbea2 */
            {8'h00}, /* 0xbea1 */
            {8'h00}, /* 0xbea0 */
            {8'h00}, /* 0xbe9f */
            {8'h00}, /* 0xbe9e */
            {8'h00}, /* 0xbe9d */
            {8'h00}, /* 0xbe9c */
            {8'h00}, /* 0xbe9b */
            {8'h00}, /* 0xbe9a */
            {8'h00}, /* 0xbe99 */
            {8'h00}, /* 0xbe98 */
            {8'h00}, /* 0xbe97 */
            {8'h00}, /* 0xbe96 */
            {8'h00}, /* 0xbe95 */
            {8'h00}, /* 0xbe94 */
            {8'h00}, /* 0xbe93 */
            {8'h00}, /* 0xbe92 */
            {8'h00}, /* 0xbe91 */
            {8'h00}, /* 0xbe90 */
            {8'h00}, /* 0xbe8f */
            {8'h00}, /* 0xbe8e */
            {8'h00}, /* 0xbe8d */
            {8'h00}, /* 0xbe8c */
            {8'h00}, /* 0xbe8b */
            {8'h00}, /* 0xbe8a */
            {8'h00}, /* 0xbe89 */
            {8'h00}, /* 0xbe88 */
            {8'h00}, /* 0xbe87 */
            {8'h00}, /* 0xbe86 */
            {8'h00}, /* 0xbe85 */
            {8'h00}, /* 0xbe84 */
            {8'h00}, /* 0xbe83 */
            {8'h00}, /* 0xbe82 */
            {8'h00}, /* 0xbe81 */
            {8'h00}, /* 0xbe80 */
            {8'h00}, /* 0xbe7f */
            {8'h00}, /* 0xbe7e */
            {8'h00}, /* 0xbe7d */
            {8'h00}, /* 0xbe7c */
            {8'h00}, /* 0xbe7b */
            {8'h00}, /* 0xbe7a */
            {8'h00}, /* 0xbe79 */
            {8'h00}, /* 0xbe78 */
            {8'h00}, /* 0xbe77 */
            {8'h00}, /* 0xbe76 */
            {8'h00}, /* 0xbe75 */
            {8'h00}, /* 0xbe74 */
            {8'h00}, /* 0xbe73 */
            {8'h00}, /* 0xbe72 */
            {8'h00}, /* 0xbe71 */
            {8'h00}, /* 0xbe70 */
            {8'h00}, /* 0xbe6f */
            {8'h00}, /* 0xbe6e */
            {8'h00}, /* 0xbe6d */
            {8'h00}, /* 0xbe6c */
            {8'h00}, /* 0xbe6b */
            {8'h00}, /* 0xbe6a */
            {8'h00}, /* 0xbe69 */
            {8'h00}, /* 0xbe68 */
            {8'h00}, /* 0xbe67 */
            {8'h00}, /* 0xbe66 */
            {8'h00}, /* 0xbe65 */
            {8'h00}, /* 0xbe64 */
            {8'h00}, /* 0xbe63 */
            {8'h00}, /* 0xbe62 */
            {8'h00}, /* 0xbe61 */
            {8'h00}, /* 0xbe60 */
            {8'h00}, /* 0xbe5f */
            {8'h00}, /* 0xbe5e */
            {8'h00}, /* 0xbe5d */
            {8'h00}, /* 0xbe5c */
            {8'h00}, /* 0xbe5b */
            {8'h00}, /* 0xbe5a */
            {8'h00}, /* 0xbe59 */
            {8'h00}, /* 0xbe58 */
            {8'h00}, /* 0xbe57 */
            {8'h00}, /* 0xbe56 */
            {8'h00}, /* 0xbe55 */
            {8'h00}, /* 0xbe54 */
            {8'h00}, /* 0xbe53 */
            {8'h00}, /* 0xbe52 */
            {8'h00}, /* 0xbe51 */
            {8'h00}, /* 0xbe50 */
            {8'h00}, /* 0xbe4f */
            {8'h00}, /* 0xbe4e */
            {8'h00}, /* 0xbe4d */
            {8'h00}, /* 0xbe4c */
            {8'h00}, /* 0xbe4b */
            {8'h00}, /* 0xbe4a */
            {8'h00}, /* 0xbe49 */
            {8'h00}, /* 0xbe48 */
            {8'h00}, /* 0xbe47 */
            {8'h00}, /* 0xbe46 */
            {8'h00}, /* 0xbe45 */
            {8'h00}, /* 0xbe44 */
            {8'h00}, /* 0xbe43 */
            {8'h00}, /* 0xbe42 */
            {8'h00}, /* 0xbe41 */
            {8'h00}, /* 0xbe40 */
            {8'h00}, /* 0xbe3f */
            {8'h00}, /* 0xbe3e */
            {8'h00}, /* 0xbe3d */
            {8'h00}, /* 0xbe3c */
            {8'h00}, /* 0xbe3b */
            {8'h00}, /* 0xbe3a */
            {8'h00}, /* 0xbe39 */
            {8'h00}, /* 0xbe38 */
            {8'h00}, /* 0xbe37 */
            {8'h00}, /* 0xbe36 */
            {8'h00}, /* 0xbe35 */
            {8'h00}, /* 0xbe34 */
            {8'h00}, /* 0xbe33 */
            {8'h00}, /* 0xbe32 */
            {8'h00}, /* 0xbe31 */
            {8'h00}, /* 0xbe30 */
            {8'h00}, /* 0xbe2f */
            {8'h00}, /* 0xbe2e */
            {8'h00}, /* 0xbe2d */
            {8'h00}, /* 0xbe2c */
            {8'h00}, /* 0xbe2b */
            {8'h00}, /* 0xbe2a */
            {8'h00}, /* 0xbe29 */
            {8'h00}, /* 0xbe28 */
            {8'h00}, /* 0xbe27 */
            {8'h00}, /* 0xbe26 */
            {8'h00}, /* 0xbe25 */
            {8'h00}, /* 0xbe24 */
            {8'h00}, /* 0xbe23 */
            {8'h00}, /* 0xbe22 */
            {8'h00}, /* 0xbe21 */
            {8'h00}, /* 0xbe20 */
            {8'h00}, /* 0xbe1f */
            {8'h00}, /* 0xbe1e */
            {8'h00}, /* 0xbe1d */
            {8'h00}, /* 0xbe1c */
            {8'h00}, /* 0xbe1b */
            {8'h00}, /* 0xbe1a */
            {8'h00}, /* 0xbe19 */
            {8'h00}, /* 0xbe18 */
            {8'h00}, /* 0xbe17 */
            {8'h00}, /* 0xbe16 */
            {8'h00}, /* 0xbe15 */
            {8'h00}, /* 0xbe14 */
            {8'h00}, /* 0xbe13 */
            {8'h00}, /* 0xbe12 */
            {8'h00}, /* 0xbe11 */
            {8'h00}, /* 0xbe10 */
            {8'h00}, /* 0xbe0f */
            {8'h00}, /* 0xbe0e */
            {8'h00}, /* 0xbe0d */
            {8'h00}, /* 0xbe0c */
            {8'h00}, /* 0xbe0b */
            {8'h00}, /* 0xbe0a */
            {8'h00}, /* 0xbe09 */
            {8'h00}, /* 0xbe08 */
            {8'h00}, /* 0xbe07 */
            {8'h00}, /* 0xbe06 */
            {8'h00}, /* 0xbe05 */
            {8'h00}, /* 0xbe04 */
            {8'h00}, /* 0xbe03 */
            {8'h00}, /* 0xbe02 */
            {8'h00}, /* 0xbe01 */
            {8'h00}, /* 0xbe00 */
            {8'h00}, /* 0xbdff */
            {8'h00}, /* 0xbdfe */
            {8'h00}, /* 0xbdfd */
            {8'h00}, /* 0xbdfc */
            {8'h00}, /* 0xbdfb */
            {8'h00}, /* 0xbdfa */
            {8'h00}, /* 0xbdf9 */
            {8'h00}, /* 0xbdf8 */
            {8'h00}, /* 0xbdf7 */
            {8'h00}, /* 0xbdf6 */
            {8'h00}, /* 0xbdf5 */
            {8'h00}, /* 0xbdf4 */
            {8'h00}, /* 0xbdf3 */
            {8'h00}, /* 0xbdf2 */
            {8'h00}, /* 0xbdf1 */
            {8'h00}, /* 0xbdf0 */
            {8'h00}, /* 0xbdef */
            {8'h00}, /* 0xbdee */
            {8'h00}, /* 0xbded */
            {8'h00}, /* 0xbdec */
            {8'h00}, /* 0xbdeb */
            {8'h00}, /* 0xbdea */
            {8'h00}, /* 0xbde9 */
            {8'h00}, /* 0xbde8 */
            {8'h00}, /* 0xbde7 */
            {8'h00}, /* 0xbde6 */
            {8'h00}, /* 0xbde5 */
            {8'h00}, /* 0xbde4 */
            {8'h00}, /* 0xbde3 */
            {8'h00}, /* 0xbde2 */
            {8'h00}, /* 0xbde1 */
            {8'h00}, /* 0xbde0 */
            {8'h00}, /* 0xbddf */
            {8'h00}, /* 0xbdde */
            {8'h00}, /* 0xbddd */
            {8'h00}, /* 0xbddc */
            {8'h00}, /* 0xbddb */
            {8'h00}, /* 0xbdda */
            {8'h00}, /* 0xbdd9 */
            {8'h00}, /* 0xbdd8 */
            {8'h00}, /* 0xbdd7 */
            {8'h00}, /* 0xbdd6 */
            {8'h00}, /* 0xbdd5 */
            {8'h00}, /* 0xbdd4 */
            {8'h00}, /* 0xbdd3 */
            {8'h00}, /* 0xbdd2 */
            {8'h00}, /* 0xbdd1 */
            {8'h00}, /* 0xbdd0 */
            {8'h00}, /* 0xbdcf */
            {8'h00}, /* 0xbdce */
            {8'h00}, /* 0xbdcd */
            {8'h00}, /* 0xbdcc */
            {8'h00}, /* 0xbdcb */
            {8'h00}, /* 0xbdca */
            {8'h00}, /* 0xbdc9 */
            {8'h00}, /* 0xbdc8 */
            {8'h00}, /* 0xbdc7 */
            {8'h00}, /* 0xbdc6 */
            {8'h00}, /* 0xbdc5 */
            {8'h00}, /* 0xbdc4 */
            {8'h00}, /* 0xbdc3 */
            {8'h00}, /* 0xbdc2 */
            {8'h00}, /* 0xbdc1 */
            {8'h00}, /* 0xbdc0 */
            {8'h00}, /* 0xbdbf */
            {8'h00}, /* 0xbdbe */
            {8'h00}, /* 0xbdbd */
            {8'h00}, /* 0xbdbc */
            {8'h00}, /* 0xbdbb */
            {8'h00}, /* 0xbdba */
            {8'h00}, /* 0xbdb9 */
            {8'h00}, /* 0xbdb8 */
            {8'h00}, /* 0xbdb7 */
            {8'h00}, /* 0xbdb6 */
            {8'h00}, /* 0xbdb5 */
            {8'h00}, /* 0xbdb4 */
            {8'h00}, /* 0xbdb3 */
            {8'h00}, /* 0xbdb2 */
            {8'h00}, /* 0xbdb1 */
            {8'h00}, /* 0xbdb0 */
            {8'h00}, /* 0xbdaf */
            {8'h00}, /* 0xbdae */
            {8'h00}, /* 0xbdad */
            {8'h00}, /* 0xbdac */
            {8'h00}, /* 0xbdab */
            {8'h00}, /* 0xbdaa */
            {8'h00}, /* 0xbda9 */
            {8'h00}, /* 0xbda8 */
            {8'h00}, /* 0xbda7 */
            {8'h00}, /* 0xbda6 */
            {8'h00}, /* 0xbda5 */
            {8'h00}, /* 0xbda4 */
            {8'h00}, /* 0xbda3 */
            {8'h00}, /* 0xbda2 */
            {8'h00}, /* 0xbda1 */
            {8'h00}, /* 0xbda0 */
            {8'h00}, /* 0xbd9f */
            {8'h00}, /* 0xbd9e */
            {8'h00}, /* 0xbd9d */
            {8'h00}, /* 0xbd9c */
            {8'h00}, /* 0xbd9b */
            {8'h00}, /* 0xbd9a */
            {8'h00}, /* 0xbd99 */
            {8'h00}, /* 0xbd98 */
            {8'h00}, /* 0xbd97 */
            {8'h00}, /* 0xbd96 */
            {8'h00}, /* 0xbd95 */
            {8'h00}, /* 0xbd94 */
            {8'h00}, /* 0xbd93 */
            {8'h00}, /* 0xbd92 */
            {8'h00}, /* 0xbd91 */
            {8'h00}, /* 0xbd90 */
            {8'h00}, /* 0xbd8f */
            {8'h00}, /* 0xbd8e */
            {8'h00}, /* 0xbd8d */
            {8'h00}, /* 0xbd8c */
            {8'h00}, /* 0xbd8b */
            {8'h00}, /* 0xbd8a */
            {8'h00}, /* 0xbd89 */
            {8'h00}, /* 0xbd88 */
            {8'h00}, /* 0xbd87 */
            {8'h00}, /* 0xbd86 */
            {8'h00}, /* 0xbd85 */
            {8'h00}, /* 0xbd84 */
            {8'h00}, /* 0xbd83 */
            {8'h00}, /* 0xbd82 */
            {8'h00}, /* 0xbd81 */
            {8'h00}, /* 0xbd80 */
            {8'h00}, /* 0xbd7f */
            {8'h00}, /* 0xbd7e */
            {8'h00}, /* 0xbd7d */
            {8'h00}, /* 0xbd7c */
            {8'h00}, /* 0xbd7b */
            {8'h00}, /* 0xbd7a */
            {8'h00}, /* 0xbd79 */
            {8'h00}, /* 0xbd78 */
            {8'h00}, /* 0xbd77 */
            {8'h00}, /* 0xbd76 */
            {8'h00}, /* 0xbd75 */
            {8'h00}, /* 0xbd74 */
            {8'h00}, /* 0xbd73 */
            {8'h00}, /* 0xbd72 */
            {8'h00}, /* 0xbd71 */
            {8'h00}, /* 0xbd70 */
            {8'h00}, /* 0xbd6f */
            {8'h00}, /* 0xbd6e */
            {8'h00}, /* 0xbd6d */
            {8'h00}, /* 0xbd6c */
            {8'h00}, /* 0xbd6b */
            {8'h00}, /* 0xbd6a */
            {8'h00}, /* 0xbd69 */
            {8'h00}, /* 0xbd68 */
            {8'h00}, /* 0xbd67 */
            {8'h00}, /* 0xbd66 */
            {8'h00}, /* 0xbd65 */
            {8'h00}, /* 0xbd64 */
            {8'h00}, /* 0xbd63 */
            {8'h00}, /* 0xbd62 */
            {8'h00}, /* 0xbd61 */
            {8'h00}, /* 0xbd60 */
            {8'h00}, /* 0xbd5f */
            {8'h00}, /* 0xbd5e */
            {8'h00}, /* 0xbd5d */
            {8'h00}, /* 0xbd5c */
            {8'h00}, /* 0xbd5b */
            {8'h00}, /* 0xbd5a */
            {8'h00}, /* 0xbd59 */
            {8'h00}, /* 0xbd58 */
            {8'h00}, /* 0xbd57 */
            {8'h00}, /* 0xbd56 */
            {8'h00}, /* 0xbd55 */
            {8'h00}, /* 0xbd54 */
            {8'h00}, /* 0xbd53 */
            {8'h00}, /* 0xbd52 */
            {8'h00}, /* 0xbd51 */
            {8'h00}, /* 0xbd50 */
            {8'h00}, /* 0xbd4f */
            {8'h00}, /* 0xbd4e */
            {8'h00}, /* 0xbd4d */
            {8'h00}, /* 0xbd4c */
            {8'h00}, /* 0xbd4b */
            {8'h00}, /* 0xbd4a */
            {8'h00}, /* 0xbd49 */
            {8'h00}, /* 0xbd48 */
            {8'h00}, /* 0xbd47 */
            {8'h00}, /* 0xbd46 */
            {8'h00}, /* 0xbd45 */
            {8'h00}, /* 0xbd44 */
            {8'h00}, /* 0xbd43 */
            {8'h00}, /* 0xbd42 */
            {8'h00}, /* 0xbd41 */
            {8'h00}, /* 0xbd40 */
            {8'h00}, /* 0xbd3f */
            {8'h00}, /* 0xbd3e */
            {8'h00}, /* 0xbd3d */
            {8'h00}, /* 0xbd3c */
            {8'h00}, /* 0xbd3b */
            {8'h00}, /* 0xbd3a */
            {8'h00}, /* 0xbd39 */
            {8'h00}, /* 0xbd38 */
            {8'h00}, /* 0xbd37 */
            {8'h00}, /* 0xbd36 */
            {8'h00}, /* 0xbd35 */
            {8'h00}, /* 0xbd34 */
            {8'h00}, /* 0xbd33 */
            {8'h00}, /* 0xbd32 */
            {8'h00}, /* 0xbd31 */
            {8'h00}, /* 0xbd30 */
            {8'h00}, /* 0xbd2f */
            {8'h00}, /* 0xbd2e */
            {8'h00}, /* 0xbd2d */
            {8'h00}, /* 0xbd2c */
            {8'h00}, /* 0xbd2b */
            {8'h00}, /* 0xbd2a */
            {8'h00}, /* 0xbd29 */
            {8'h00}, /* 0xbd28 */
            {8'h00}, /* 0xbd27 */
            {8'h00}, /* 0xbd26 */
            {8'h00}, /* 0xbd25 */
            {8'h00}, /* 0xbd24 */
            {8'h00}, /* 0xbd23 */
            {8'h00}, /* 0xbd22 */
            {8'h00}, /* 0xbd21 */
            {8'h00}, /* 0xbd20 */
            {8'h00}, /* 0xbd1f */
            {8'h00}, /* 0xbd1e */
            {8'h00}, /* 0xbd1d */
            {8'h00}, /* 0xbd1c */
            {8'h00}, /* 0xbd1b */
            {8'h00}, /* 0xbd1a */
            {8'h00}, /* 0xbd19 */
            {8'h00}, /* 0xbd18 */
            {8'h00}, /* 0xbd17 */
            {8'h00}, /* 0xbd16 */
            {8'h00}, /* 0xbd15 */
            {8'h00}, /* 0xbd14 */
            {8'h00}, /* 0xbd13 */
            {8'h00}, /* 0xbd12 */
            {8'h00}, /* 0xbd11 */
            {8'h00}, /* 0xbd10 */
            {8'h00}, /* 0xbd0f */
            {8'h00}, /* 0xbd0e */
            {8'h00}, /* 0xbd0d */
            {8'h00}, /* 0xbd0c */
            {8'h00}, /* 0xbd0b */
            {8'h00}, /* 0xbd0a */
            {8'h00}, /* 0xbd09 */
            {8'h00}, /* 0xbd08 */
            {8'h00}, /* 0xbd07 */
            {8'h00}, /* 0xbd06 */
            {8'h00}, /* 0xbd05 */
            {8'h00}, /* 0xbd04 */
            {8'h00}, /* 0xbd03 */
            {8'h00}, /* 0xbd02 */
            {8'h00}, /* 0xbd01 */
            {8'h00}, /* 0xbd00 */
            {8'h00}, /* 0xbcff */
            {8'h00}, /* 0xbcfe */
            {8'h00}, /* 0xbcfd */
            {8'h00}, /* 0xbcfc */
            {8'h00}, /* 0xbcfb */
            {8'h00}, /* 0xbcfa */
            {8'h00}, /* 0xbcf9 */
            {8'h00}, /* 0xbcf8 */
            {8'h00}, /* 0xbcf7 */
            {8'h00}, /* 0xbcf6 */
            {8'h00}, /* 0xbcf5 */
            {8'h00}, /* 0xbcf4 */
            {8'h00}, /* 0xbcf3 */
            {8'h00}, /* 0xbcf2 */
            {8'h00}, /* 0xbcf1 */
            {8'h00}, /* 0xbcf0 */
            {8'h00}, /* 0xbcef */
            {8'h00}, /* 0xbcee */
            {8'h00}, /* 0xbced */
            {8'h00}, /* 0xbcec */
            {8'h00}, /* 0xbceb */
            {8'h00}, /* 0xbcea */
            {8'h00}, /* 0xbce9 */
            {8'h00}, /* 0xbce8 */
            {8'h00}, /* 0xbce7 */
            {8'h00}, /* 0xbce6 */
            {8'h00}, /* 0xbce5 */
            {8'h00}, /* 0xbce4 */
            {8'h00}, /* 0xbce3 */
            {8'h00}, /* 0xbce2 */
            {8'h00}, /* 0xbce1 */
            {8'h00}, /* 0xbce0 */
            {8'h00}, /* 0xbcdf */
            {8'h00}, /* 0xbcde */
            {8'h00}, /* 0xbcdd */
            {8'h00}, /* 0xbcdc */
            {8'h00}, /* 0xbcdb */
            {8'h00}, /* 0xbcda */
            {8'h00}, /* 0xbcd9 */
            {8'h00}, /* 0xbcd8 */
            {8'h00}, /* 0xbcd7 */
            {8'h00}, /* 0xbcd6 */
            {8'h00}, /* 0xbcd5 */
            {8'h00}, /* 0xbcd4 */
            {8'h00}, /* 0xbcd3 */
            {8'h00}, /* 0xbcd2 */
            {8'h00}, /* 0xbcd1 */
            {8'h00}, /* 0xbcd0 */
            {8'h00}, /* 0xbccf */
            {8'h00}, /* 0xbcce */
            {8'h00}, /* 0xbccd */
            {8'h00}, /* 0xbccc */
            {8'h00}, /* 0xbccb */
            {8'h00}, /* 0xbcca */
            {8'h00}, /* 0xbcc9 */
            {8'h00}, /* 0xbcc8 */
            {8'h00}, /* 0xbcc7 */
            {8'h00}, /* 0xbcc6 */
            {8'h00}, /* 0xbcc5 */
            {8'h00}, /* 0xbcc4 */
            {8'h00}, /* 0xbcc3 */
            {8'h00}, /* 0xbcc2 */
            {8'h00}, /* 0xbcc1 */
            {8'h00}, /* 0xbcc0 */
            {8'h00}, /* 0xbcbf */
            {8'h00}, /* 0xbcbe */
            {8'h00}, /* 0xbcbd */
            {8'h00}, /* 0xbcbc */
            {8'h00}, /* 0xbcbb */
            {8'h00}, /* 0xbcba */
            {8'h00}, /* 0xbcb9 */
            {8'h00}, /* 0xbcb8 */
            {8'h00}, /* 0xbcb7 */
            {8'h00}, /* 0xbcb6 */
            {8'h00}, /* 0xbcb5 */
            {8'h00}, /* 0xbcb4 */
            {8'h00}, /* 0xbcb3 */
            {8'h00}, /* 0xbcb2 */
            {8'h00}, /* 0xbcb1 */
            {8'h00}, /* 0xbcb0 */
            {8'h00}, /* 0xbcaf */
            {8'h00}, /* 0xbcae */
            {8'h00}, /* 0xbcad */
            {8'h00}, /* 0xbcac */
            {8'h00}, /* 0xbcab */
            {8'h00}, /* 0xbcaa */
            {8'h00}, /* 0xbca9 */
            {8'h00}, /* 0xbca8 */
            {8'h00}, /* 0xbca7 */
            {8'h00}, /* 0xbca6 */
            {8'h00}, /* 0xbca5 */
            {8'h00}, /* 0xbca4 */
            {8'h00}, /* 0xbca3 */
            {8'h00}, /* 0xbca2 */
            {8'h00}, /* 0xbca1 */
            {8'h00}, /* 0xbca0 */
            {8'h00}, /* 0xbc9f */
            {8'h00}, /* 0xbc9e */
            {8'h00}, /* 0xbc9d */
            {8'h00}, /* 0xbc9c */
            {8'h00}, /* 0xbc9b */
            {8'h00}, /* 0xbc9a */
            {8'h00}, /* 0xbc99 */
            {8'h00}, /* 0xbc98 */
            {8'h00}, /* 0xbc97 */
            {8'h00}, /* 0xbc96 */
            {8'h00}, /* 0xbc95 */
            {8'h00}, /* 0xbc94 */
            {8'h00}, /* 0xbc93 */
            {8'h00}, /* 0xbc92 */
            {8'h00}, /* 0xbc91 */
            {8'h00}, /* 0xbc90 */
            {8'h00}, /* 0xbc8f */
            {8'h00}, /* 0xbc8e */
            {8'h00}, /* 0xbc8d */
            {8'h00}, /* 0xbc8c */
            {8'h00}, /* 0xbc8b */
            {8'h00}, /* 0xbc8a */
            {8'h00}, /* 0xbc89 */
            {8'h00}, /* 0xbc88 */
            {8'h00}, /* 0xbc87 */
            {8'h00}, /* 0xbc86 */
            {8'h00}, /* 0xbc85 */
            {8'h00}, /* 0xbc84 */
            {8'h00}, /* 0xbc83 */
            {8'h00}, /* 0xbc82 */
            {8'h00}, /* 0xbc81 */
            {8'h00}, /* 0xbc80 */
            {8'h00}, /* 0xbc7f */
            {8'h00}, /* 0xbc7e */
            {8'h00}, /* 0xbc7d */
            {8'h00}, /* 0xbc7c */
            {8'h00}, /* 0xbc7b */
            {8'h00}, /* 0xbc7a */
            {8'h00}, /* 0xbc79 */
            {8'h00}, /* 0xbc78 */
            {8'h00}, /* 0xbc77 */
            {8'h00}, /* 0xbc76 */
            {8'h00}, /* 0xbc75 */
            {8'h00}, /* 0xbc74 */
            {8'h00}, /* 0xbc73 */
            {8'h00}, /* 0xbc72 */
            {8'h00}, /* 0xbc71 */
            {8'h00}, /* 0xbc70 */
            {8'h00}, /* 0xbc6f */
            {8'h00}, /* 0xbc6e */
            {8'h00}, /* 0xbc6d */
            {8'h00}, /* 0xbc6c */
            {8'h00}, /* 0xbc6b */
            {8'h00}, /* 0xbc6a */
            {8'h00}, /* 0xbc69 */
            {8'h00}, /* 0xbc68 */
            {8'h00}, /* 0xbc67 */
            {8'h00}, /* 0xbc66 */
            {8'h00}, /* 0xbc65 */
            {8'h00}, /* 0xbc64 */
            {8'h00}, /* 0xbc63 */
            {8'h00}, /* 0xbc62 */
            {8'h00}, /* 0xbc61 */
            {8'h00}, /* 0xbc60 */
            {8'h00}, /* 0xbc5f */
            {8'h00}, /* 0xbc5e */
            {8'h00}, /* 0xbc5d */
            {8'h00}, /* 0xbc5c */
            {8'h00}, /* 0xbc5b */
            {8'h00}, /* 0xbc5a */
            {8'h00}, /* 0xbc59 */
            {8'h00}, /* 0xbc58 */
            {8'h00}, /* 0xbc57 */
            {8'h00}, /* 0xbc56 */
            {8'h00}, /* 0xbc55 */
            {8'h00}, /* 0xbc54 */
            {8'h00}, /* 0xbc53 */
            {8'h00}, /* 0xbc52 */
            {8'h00}, /* 0xbc51 */
            {8'h00}, /* 0xbc50 */
            {8'h00}, /* 0xbc4f */
            {8'h00}, /* 0xbc4e */
            {8'h00}, /* 0xbc4d */
            {8'h00}, /* 0xbc4c */
            {8'h00}, /* 0xbc4b */
            {8'h00}, /* 0xbc4a */
            {8'h00}, /* 0xbc49 */
            {8'h00}, /* 0xbc48 */
            {8'h00}, /* 0xbc47 */
            {8'h00}, /* 0xbc46 */
            {8'h00}, /* 0xbc45 */
            {8'h00}, /* 0xbc44 */
            {8'h00}, /* 0xbc43 */
            {8'h00}, /* 0xbc42 */
            {8'h00}, /* 0xbc41 */
            {8'h00}, /* 0xbc40 */
            {8'h00}, /* 0xbc3f */
            {8'h00}, /* 0xbc3e */
            {8'h00}, /* 0xbc3d */
            {8'h00}, /* 0xbc3c */
            {8'h00}, /* 0xbc3b */
            {8'h00}, /* 0xbc3a */
            {8'h00}, /* 0xbc39 */
            {8'h00}, /* 0xbc38 */
            {8'h00}, /* 0xbc37 */
            {8'h00}, /* 0xbc36 */
            {8'h00}, /* 0xbc35 */
            {8'h00}, /* 0xbc34 */
            {8'h00}, /* 0xbc33 */
            {8'h00}, /* 0xbc32 */
            {8'h00}, /* 0xbc31 */
            {8'h00}, /* 0xbc30 */
            {8'h00}, /* 0xbc2f */
            {8'h00}, /* 0xbc2e */
            {8'h00}, /* 0xbc2d */
            {8'h00}, /* 0xbc2c */
            {8'h00}, /* 0xbc2b */
            {8'h00}, /* 0xbc2a */
            {8'h00}, /* 0xbc29 */
            {8'h00}, /* 0xbc28 */
            {8'h00}, /* 0xbc27 */
            {8'h00}, /* 0xbc26 */
            {8'h00}, /* 0xbc25 */
            {8'h00}, /* 0xbc24 */
            {8'h00}, /* 0xbc23 */
            {8'h00}, /* 0xbc22 */
            {8'h00}, /* 0xbc21 */
            {8'h00}, /* 0xbc20 */
            {8'h00}, /* 0xbc1f */
            {8'h00}, /* 0xbc1e */
            {8'h00}, /* 0xbc1d */
            {8'h00}, /* 0xbc1c */
            {8'h00}, /* 0xbc1b */
            {8'h00}, /* 0xbc1a */
            {8'h00}, /* 0xbc19 */
            {8'h00}, /* 0xbc18 */
            {8'h00}, /* 0xbc17 */
            {8'h00}, /* 0xbc16 */
            {8'h00}, /* 0xbc15 */
            {8'h00}, /* 0xbc14 */
            {8'h00}, /* 0xbc13 */
            {8'h00}, /* 0xbc12 */
            {8'h00}, /* 0xbc11 */
            {8'h00}, /* 0xbc10 */
            {8'h00}, /* 0xbc0f */
            {8'h00}, /* 0xbc0e */
            {8'h00}, /* 0xbc0d */
            {8'h00}, /* 0xbc0c */
            {8'h00}, /* 0xbc0b */
            {8'h00}, /* 0xbc0a */
            {8'h00}, /* 0xbc09 */
            {8'h00}, /* 0xbc08 */
            {8'h00}, /* 0xbc07 */
            {8'h00}, /* 0xbc06 */
            {8'h00}, /* 0xbc05 */
            {8'h00}, /* 0xbc04 */
            {8'h00}, /* 0xbc03 */
            {8'h00}, /* 0xbc02 */
            {8'h00}, /* 0xbc01 */
            {8'h00}, /* 0xbc00 */
            {8'h00}, /* 0xbbff */
            {8'h00}, /* 0xbbfe */
            {8'h00}, /* 0xbbfd */
            {8'h00}, /* 0xbbfc */
            {8'h00}, /* 0xbbfb */
            {8'h00}, /* 0xbbfa */
            {8'h00}, /* 0xbbf9 */
            {8'h00}, /* 0xbbf8 */
            {8'h00}, /* 0xbbf7 */
            {8'h00}, /* 0xbbf6 */
            {8'h00}, /* 0xbbf5 */
            {8'h00}, /* 0xbbf4 */
            {8'h00}, /* 0xbbf3 */
            {8'h00}, /* 0xbbf2 */
            {8'h00}, /* 0xbbf1 */
            {8'h00}, /* 0xbbf0 */
            {8'h00}, /* 0xbbef */
            {8'h00}, /* 0xbbee */
            {8'h00}, /* 0xbbed */
            {8'h00}, /* 0xbbec */
            {8'h00}, /* 0xbbeb */
            {8'h00}, /* 0xbbea */
            {8'h00}, /* 0xbbe9 */
            {8'h00}, /* 0xbbe8 */
            {8'h00}, /* 0xbbe7 */
            {8'h00}, /* 0xbbe6 */
            {8'h00}, /* 0xbbe5 */
            {8'h00}, /* 0xbbe4 */
            {8'h00}, /* 0xbbe3 */
            {8'h00}, /* 0xbbe2 */
            {8'h00}, /* 0xbbe1 */
            {8'h00}, /* 0xbbe0 */
            {8'h00}, /* 0xbbdf */
            {8'h00}, /* 0xbbde */
            {8'h00}, /* 0xbbdd */
            {8'h00}, /* 0xbbdc */
            {8'h00}, /* 0xbbdb */
            {8'h00}, /* 0xbbda */
            {8'h00}, /* 0xbbd9 */
            {8'h00}, /* 0xbbd8 */
            {8'h00}, /* 0xbbd7 */
            {8'h00}, /* 0xbbd6 */
            {8'h00}, /* 0xbbd5 */
            {8'h00}, /* 0xbbd4 */
            {8'h00}, /* 0xbbd3 */
            {8'h00}, /* 0xbbd2 */
            {8'h00}, /* 0xbbd1 */
            {8'h00}, /* 0xbbd0 */
            {8'h00}, /* 0xbbcf */
            {8'h00}, /* 0xbbce */
            {8'h00}, /* 0xbbcd */
            {8'h00}, /* 0xbbcc */
            {8'h00}, /* 0xbbcb */
            {8'h00}, /* 0xbbca */
            {8'h00}, /* 0xbbc9 */
            {8'h00}, /* 0xbbc8 */
            {8'h00}, /* 0xbbc7 */
            {8'h00}, /* 0xbbc6 */
            {8'h00}, /* 0xbbc5 */
            {8'h00}, /* 0xbbc4 */
            {8'h00}, /* 0xbbc3 */
            {8'h00}, /* 0xbbc2 */
            {8'h00}, /* 0xbbc1 */
            {8'h00}, /* 0xbbc0 */
            {8'h00}, /* 0xbbbf */
            {8'h00}, /* 0xbbbe */
            {8'h00}, /* 0xbbbd */
            {8'h00}, /* 0xbbbc */
            {8'h00}, /* 0xbbbb */
            {8'h00}, /* 0xbbba */
            {8'h00}, /* 0xbbb9 */
            {8'h00}, /* 0xbbb8 */
            {8'h00}, /* 0xbbb7 */
            {8'h00}, /* 0xbbb6 */
            {8'h00}, /* 0xbbb5 */
            {8'h00}, /* 0xbbb4 */
            {8'h00}, /* 0xbbb3 */
            {8'h00}, /* 0xbbb2 */
            {8'h00}, /* 0xbbb1 */
            {8'h00}, /* 0xbbb0 */
            {8'h00}, /* 0xbbaf */
            {8'h00}, /* 0xbbae */
            {8'h00}, /* 0xbbad */
            {8'h00}, /* 0xbbac */
            {8'h00}, /* 0xbbab */
            {8'h00}, /* 0xbbaa */
            {8'h00}, /* 0xbba9 */
            {8'h00}, /* 0xbba8 */
            {8'h00}, /* 0xbba7 */
            {8'h00}, /* 0xbba6 */
            {8'h00}, /* 0xbba5 */
            {8'h00}, /* 0xbba4 */
            {8'h00}, /* 0xbba3 */
            {8'h00}, /* 0xbba2 */
            {8'h00}, /* 0xbba1 */
            {8'h00}, /* 0xbba0 */
            {8'h00}, /* 0xbb9f */
            {8'h00}, /* 0xbb9e */
            {8'h00}, /* 0xbb9d */
            {8'h00}, /* 0xbb9c */
            {8'h00}, /* 0xbb9b */
            {8'h00}, /* 0xbb9a */
            {8'h00}, /* 0xbb99 */
            {8'h00}, /* 0xbb98 */
            {8'h00}, /* 0xbb97 */
            {8'h00}, /* 0xbb96 */
            {8'h00}, /* 0xbb95 */
            {8'h00}, /* 0xbb94 */
            {8'h00}, /* 0xbb93 */
            {8'h00}, /* 0xbb92 */
            {8'h00}, /* 0xbb91 */
            {8'h00}, /* 0xbb90 */
            {8'h00}, /* 0xbb8f */
            {8'h00}, /* 0xbb8e */
            {8'h00}, /* 0xbb8d */
            {8'h00}, /* 0xbb8c */
            {8'h00}, /* 0xbb8b */
            {8'h00}, /* 0xbb8a */
            {8'h00}, /* 0xbb89 */
            {8'h00}, /* 0xbb88 */
            {8'h00}, /* 0xbb87 */
            {8'h00}, /* 0xbb86 */
            {8'h00}, /* 0xbb85 */
            {8'h00}, /* 0xbb84 */
            {8'h00}, /* 0xbb83 */
            {8'h00}, /* 0xbb82 */
            {8'h00}, /* 0xbb81 */
            {8'h00}, /* 0xbb80 */
            {8'h00}, /* 0xbb7f */
            {8'h00}, /* 0xbb7e */
            {8'h00}, /* 0xbb7d */
            {8'h00}, /* 0xbb7c */
            {8'h00}, /* 0xbb7b */
            {8'h00}, /* 0xbb7a */
            {8'h00}, /* 0xbb79 */
            {8'h00}, /* 0xbb78 */
            {8'h00}, /* 0xbb77 */
            {8'h00}, /* 0xbb76 */
            {8'h00}, /* 0xbb75 */
            {8'h00}, /* 0xbb74 */
            {8'h00}, /* 0xbb73 */
            {8'h00}, /* 0xbb72 */
            {8'h00}, /* 0xbb71 */
            {8'h00}, /* 0xbb70 */
            {8'h00}, /* 0xbb6f */
            {8'h00}, /* 0xbb6e */
            {8'h00}, /* 0xbb6d */
            {8'h00}, /* 0xbb6c */
            {8'h00}, /* 0xbb6b */
            {8'h00}, /* 0xbb6a */
            {8'h00}, /* 0xbb69 */
            {8'h00}, /* 0xbb68 */
            {8'h00}, /* 0xbb67 */
            {8'h00}, /* 0xbb66 */
            {8'h00}, /* 0xbb65 */
            {8'h00}, /* 0xbb64 */
            {8'h00}, /* 0xbb63 */
            {8'h00}, /* 0xbb62 */
            {8'h00}, /* 0xbb61 */
            {8'h00}, /* 0xbb60 */
            {8'h00}, /* 0xbb5f */
            {8'h00}, /* 0xbb5e */
            {8'h00}, /* 0xbb5d */
            {8'h00}, /* 0xbb5c */
            {8'h00}, /* 0xbb5b */
            {8'h00}, /* 0xbb5a */
            {8'h00}, /* 0xbb59 */
            {8'h00}, /* 0xbb58 */
            {8'h00}, /* 0xbb57 */
            {8'h00}, /* 0xbb56 */
            {8'h00}, /* 0xbb55 */
            {8'h00}, /* 0xbb54 */
            {8'h00}, /* 0xbb53 */
            {8'h00}, /* 0xbb52 */
            {8'h00}, /* 0xbb51 */
            {8'h00}, /* 0xbb50 */
            {8'h00}, /* 0xbb4f */
            {8'h00}, /* 0xbb4e */
            {8'h00}, /* 0xbb4d */
            {8'h00}, /* 0xbb4c */
            {8'h00}, /* 0xbb4b */
            {8'h00}, /* 0xbb4a */
            {8'h00}, /* 0xbb49 */
            {8'h00}, /* 0xbb48 */
            {8'h00}, /* 0xbb47 */
            {8'h00}, /* 0xbb46 */
            {8'h00}, /* 0xbb45 */
            {8'h00}, /* 0xbb44 */
            {8'h00}, /* 0xbb43 */
            {8'h00}, /* 0xbb42 */
            {8'h00}, /* 0xbb41 */
            {8'h00}, /* 0xbb40 */
            {8'h00}, /* 0xbb3f */
            {8'h00}, /* 0xbb3e */
            {8'h00}, /* 0xbb3d */
            {8'h00}, /* 0xbb3c */
            {8'h00}, /* 0xbb3b */
            {8'h00}, /* 0xbb3a */
            {8'h00}, /* 0xbb39 */
            {8'h00}, /* 0xbb38 */
            {8'h00}, /* 0xbb37 */
            {8'h00}, /* 0xbb36 */
            {8'h00}, /* 0xbb35 */
            {8'h00}, /* 0xbb34 */
            {8'h00}, /* 0xbb33 */
            {8'h00}, /* 0xbb32 */
            {8'h00}, /* 0xbb31 */
            {8'h00}, /* 0xbb30 */
            {8'h00}, /* 0xbb2f */
            {8'h00}, /* 0xbb2e */
            {8'h00}, /* 0xbb2d */
            {8'h00}, /* 0xbb2c */
            {8'h00}, /* 0xbb2b */
            {8'h00}, /* 0xbb2a */
            {8'h00}, /* 0xbb29 */
            {8'h00}, /* 0xbb28 */
            {8'h00}, /* 0xbb27 */
            {8'h00}, /* 0xbb26 */
            {8'h00}, /* 0xbb25 */
            {8'h00}, /* 0xbb24 */
            {8'h00}, /* 0xbb23 */
            {8'h00}, /* 0xbb22 */
            {8'h00}, /* 0xbb21 */
            {8'h00}, /* 0xbb20 */
            {8'h00}, /* 0xbb1f */
            {8'h00}, /* 0xbb1e */
            {8'h00}, /* 0xbb1d */
            {8'h00}, /* 0xbb1c */
            {8'h00}, /* 0xbb1b */
            {8'h00}, /* 0xbb1a */
            {8'h00}, /* 0xbb19 */
            {8'h00}, /* 0xbb18 */
            {8'h00}, /* 0xbb17 */
            {8'h00}, /* 0xbb16 */
            {8'h00}, /* 0xbb15 */
            {8'h00}, /* 0xbb14 */
            {8'h00}, /* 0xbb13 */
            {8'h00}, /* 0xbb12 */
            {8'h00}, /* 0xbb11 */
            {8'h00}, /* 0xbb10 */
            {8'h00}, /* 0xbb0f */
            {8'h00}, /* 0xbb0e */
            {8'h00}, /* 0xbb0d */
            {8'h00}, /* 0xbb0c */
            {8'h00}, /* 0xbb0b */
            {8'h00}, /* 0xbb0a */
            {8'h00}, /* 0xbb09 */
            {8'h00}, /* 0xbb08 */
            {8'h00}, /* 0xbb07 */
            {8'h00}, /* 0xbb06 */
            {8'h00}, /* 0xbb05 */
            {8'h00}, /* 0xbb04 */
            {8'h00}, /* 0xbb03 */
            {8'h00}, /* 0xbb02 */
            {8'h00}, /* 0xbb01 */
            {8'h00}, /* 0xbb00 */
            {8'h00}, /* 0xbaff */
            {8'h00}, /* 0xbafe */
            {8'h00}, /* 0xbafd */
            {8'h00}, /* 0xbafc */
            {8'h00}, /* 0xbafb */
            {8'h00}, /* 0xbafa */
            {8'h00}, /* 0xbaf9 */
            {8'h00}, /* 0xbaf8 */
            {8'h00}, /* 0xbaf7 */
            {8'h00}, /* 0xbaf6 */
            {8'h00}, /* 0xbaf5 */
            {8'h00}, /* 0xbaf4 */
            {8'h00}, /* 0xbaf3 */
            {8'h00}, /* 0xbaf2 */
            {8'h00}, /* 0xbaf1 */
            {8'h00}, /* 0xbaf0 */
            {8'h00}, /* 0xbaef */
            {8'h00}, /* 0xbaee */
            {8'h00}, /* 0xbaed */
            {8'h00}, /* 0xbaec */
            {8'h00}, /* 0xbaeb */
            {8'h00}, /* 0xbaea */
            {8'h00}, /* 0xbae9 */
            {8'h00}, /* 0xbae8 */
            {8'h00}, /* 0xbae7 */
            {8'h00}, /* 0xbae6 */
            {8'h00}, /* 0xbae5 */
            {8'h00}, /* 0xbae4 */
            {8'h00}, /* 0xbae3 */
            {8'h00}, /* 0xbae2 */
            {8'h00}, /* 0xbae1 */
            {8'h00}, /* 0xbae0 */
            {8'h00}, /* 0xbadf */
            {8'h00}, /* 0xbade */
            {8'h00}, /* 0xbadd */
            {8'h00}, /* 0xbadc */
            {8'h00}, /* 0xbadb */
            {8'h00}, /* 0xbada */
            {8'h00}, /* 0xbad9 */
            {8'h00}, /* 0xbad8 */
            {8'h00}, /* 0xbad7 */
            {8'h00}, /* 0xbad6 */
            {8'h00}, /* 0xbad5 */
            {8'h00}, /* 0xbad4 */
            {8'h00}, /* 0xbad3 */
            {8'h00}, /* 0xbad2 */
            {8'h00}, /* 0xbad1 */
            {8'h00}, /* 0xbad0 */
            {8'h00}, /* 0xbacf */
            {8'h00}, /* 0xbace */
            {8'h00}, /* 0xbacd */
            {8'h00}, /* 0xbacc */
            {8'h00}, /* 0xbacb */
            {8'h00}, /* 0xbaca */
            {8'h00}, /* 0xbac9 */
            {8'h00}, /* 0xbac8 */
            {8'h00}, /* 0xbac7 */
            {8'h00}, /* 0xbac6 */
            {8'h00}, /* 0xbac5 */
            {8'h00}, /* 0xbac4 */
            {8'h00}, /* 0xbac3 */
            {8'h00}, /* 0xbac2 */
            {8'h00}, /* 0xbac1 */
            {8'h00}, /* 0xbac0 */
            {8'h00}, /* 0xbabf */
            {8'h00}, /* 0xbabe */
            {8'h00}, /* 0xbabd */
            {8'h00}, /* 0xbabc */
            {8'h00}, /* 0xbabb */
            {8'h00}, /* 0xbaba */
            {8'h00}, /* 0xbab9 */
            {8'h00}, /* 0xbab8 */
            {8'h00}, /* 0xbab7 */
            {8'h00}, /* 0xbab6 */
            {8'h00}, /* 0xbab5 */
            {8'h00}, /* 0xbab4 */
            {8'h00}, /* 0xbab3 */
            {8'h00}, /* 0xbab2 */
            {8'h00}, /* 0xbab1 */
            {8'h00}, /* 0xbab0 */
            {8'h00}, /* 0xbaaf */
            {8'h00}, /* 0xbaae */
            {8'h00}, /* 0xbaad */
            {8'h00}, /* 0xbaac */
            {8'h00}, /* 0xbaab */
            {8'h00}, /* 0xbaaa */
            {8'h00}, /* 0xbaa9 */
            {8'h00}, /* 0xbaa8 */
            {8'h00}, /* 0xbaa7 */
            {8'h00}, /* 0xbaa6 */
            {8'h00}, /* 0xbaa5 */
            {8'h00}, /* 0xbaa4 */
            {8'h00}, /* 0xbaa3 */
            {8'h00}, /* 0xbaa2 */
            {8'h00}, /* 0xbaa1 */
            {8'h00}, /* 0xbaa0 */
            {8'h00}, /* 0xba9f */
            {8'h00}, /* 0xba9e */
            {8'h00}, /* 0xba9d */
            {8'h00}, /* 0xba9c */
            {8'h00}, /* 0xba9b */
            {8'h00}, /* 0xba9a */
            {8'h00}, /* 0xba99 */
            {8'h00}, /* 0xba98 */
            {8'h00}, /* 0xba97 */
            {8'h00}, /* 0xba96 */
            {8'h00}, /* 0xba95 */
            {8'h00}, /* 0xba94 */
            {8'h00}, /* 0xba93 */
            {8'h00}, /* 0xba92 */
            {8'h00}, /* 0xba91 */
            {8'h00}, /* 0xba90 */
            {8'h00}, /* 0xba8f */
            {8'h00}, /* 0xba8e */
            {8'h00}, /* 0xba8d */
            {8'h00}, /* 0xba8c */
            {8'h00}, /* 0xba8b */
            {8'h00}, /* 0xba8a */
            {8'h00}, /* 0xba89 */
            {8'h00}, /* 0xba88 */
            {8'h00}, /* 0xba87 */
            {8'h00}, /* 0xba86 */
            {8'h00}, /* 0xba85 */
            {8'h00}, /* 0xba84 */
            {8'h00}, /* 0xba83 */
            {8'h00}, /* 0xba82 */
            {8'h00}, /* 0xba81 */
            {8'h00}, /* 0xba80 */
            {8'h00}, /* 0xba7f */
            {8'h00}, /* 0xba7e */
            {8'h00}, /* 0xba7d */
            {8'h00}, /* 0xba7c */
            {8'h00}, /* 0xba7b */
            {8'h00}, /* 0xba7a */
            {8'h00}, /* 0xba79 */
            {8'h00}, /* 0xba78 */
            {8'h00}, /* 0xba77 */
            {8'h00}, /* 0xba76 */
            {8'h00}, /* 0xba75 */
            {8'h00}, /* 0xba74 */
            {8'h00}, /* 0xba73 */
            {8'h00}, /* 0xba72 */
            {8'h00}, /* 0xba71 */
            {8'h00}, /* 0xba70 */
            {8'h00}, /* 0xba6f */
            {8'h00}, /* 0xba6e */
            {8'h00}, /* 0xba6d */
            {8'h00}, /* 0xba6c */
            {8'h00}, /* 0xba6b */
            {8'h00}, /* 0xba6a */
            {8'h00}, /* 0xba69 */
            {8'h00}, /* 0xba68 */
            {8'h00}, /* 0xba67 */
            {8'h00}, /* 0xba66 */
            {8'h00}, /* 0xba65 */
            {8'h00}, /* 0xba64 */
            {8'h00}, /* 0xba63 */
            {8'h00}, /* 0xba62 */
            {8'h00}, /* 0xba61 */
            {8'h00}, /* 0xba60 */
            {8'h00}, /* 0xba5f */
            {8'h00}, /* 0xba5e */
            {8'h00}, /* 0xba5d */
            {8'h00}, /* 0xba5c */
            {8'h00}, /* 0xba5b */
            {8'h00}, /* 0xba5a */
            {8'h00}, /* 0xba59 */
            {8'h00}, /* 0xba58 */
            {8'h00}, /* 0xba57 */
            {8'h00}, /* 0xba56 */
            {8'h00}, /* 0xba55 */
            {8'h00}, /* 0xba54 */
            {8'h00}, /* 0xba53 */
            {8'h00}, /* 0xba52 */
            {8'h00}, /* 0xba51 */
            {8'h00}, /* 0xba50 */
            {8'h00}, /* 0xba4f */
            {8'h00}, /* 0xba4e */
            {8'h00}, /* 0xba4d */
            {8'h00}, /* 0xba4c */
            {8'h00}, /* 0xba4b */
            {8'h00}, /* 0xba4a */
            {8'h00}, /* 0xba49 */
            {8'h00}, /* 0xba48 */
            {8'h00}, /* 0xba47 */
            {8'h00}, /* 0xba46 */
            {8'h00}, /* 0xba45 */
            {8'h00}, /* 0xba44 */
            {8'h00}, /* 0xba43 */
            {8'h00}, /* 0xba42 */
            {8'h00}, /* 0xba41 */
            {8'h00}, /* 0xba40 */
            {8'h00}, /* 0xba3f */
            {8'h00}, /* 0xba3e */
            {8'h00}, /* 0xba3d */
            {8'h00}, /* 0xba3c */
            {8'h00}, /* 0xba3b */
            {8'h00}, /* 0xba3a */
            {8'h00}, /* 0xba39 */
            {8'h00}, /* 0xba38 */
            {8'h00}, /* 0xba37 */
            {8'h00}, /* 0xba36 */
            {8'h00}, /* 0xba35 */
            {8'h00}, /* 0xba34 */
            {8'h00}, /* 0xba33 */
            {8'h00}, /* 0xba32 */
            {8'h00}, /* 0xba31 */
            {8'h00}, /* 0xba30 */
            {8'h00}, /* 0xba2f */
            {8'h00}, /* 0xba2e */
            {8'h00}, /* 0xba2d */
            {8'h00}, /* 0xba2c */
            {8'h00}, /* 0xba2b */
            {8'h00}, /* 0xba2a */
            {8'h00}, /* 0xba29 */
            {8'h00}, /* 0xba28 */
            {8'h00}, /* 0xba27 */
            {8'h00}, /* 0xba26 */
            {8'h00}, /* 0xba25 */
            {8'h00}, /* 0xba24 */
            {8'h00}, /* 0xba23 */
            {8'h00}, /* 0xba22 */
            {8'h00}, /* 0xba21 */
            {8'h00}, /* 0xba20 */
            {8'h00}, /* 0xba1f */
            {8'h00}, /* 0xba1e */
            {8'h00}, /* 0xba1d */
            {8'h00}, /* 0xba1c */
            {8'h00}, /* 0xba1b */
            {8'h00}, /* 0xba1a */
            {8'h00}, /* 0xba19 */
            {8'h00}, /* 0xba18 */
            {8'h00}, /* 0xba17 */
            {8'h00}, /* 0xba16 */
            {8'h00}, /* 0xba15 */
            {8'h00}, /* 0xba14 */
            {8'h00}, /* 0xba13 */
            {8'h00}, /* 0xba12 */
            {8'h00}, /* 0xba11 */
            {8'h00}, /* 0xba10 */
            {8'h00}, /* 0xba0f */
            {8'h00}, /* 0xba0e */
            {8'h00}, /* 0xba0d */
            {8'h00}, /* 0xba0c */
            {8'h00}, /* 0xba0b */
            {8'h00}, /* 0xba0a */
            {8'h00}, /* 0xba09 */
            {8'h00}, /* 0xba08 */
            {8'h00}, /* 0xba07 */
            {8'h00}, /* 0xba06 */
            {8'h00}, /* 0xba05 */
            {8'h00}, /* 0xba04 */
            {8'h00}, /* 0xba03 */
            {8'h00}, /* 0xba02 */
            {8'h00}, /* 0xba01 */
            {8'h00}, /* 0xba00 */
            {8'h00}, /* 0xb9ff */
            {8'h00}, /* 0xb9fe */
            {8'h00}, /* 0xb9fd */
            {8'h00}, /* 0xb9fc */
            {8'h00}, /* 0xb9fb */
            {8'h00}, /* 0xb9fa */
            {8'h00}, /* 0xb9f9 */
            {8'h00}, /* 0xb9f8 */
            {8'h00}, /* 0xb9f7 */
            {8'h00}, /* 0xb9f6 */
            {8'h00}, /* 0xb9f5 */
            {8'h00}, /* 0xb9f4 */
            {8'h00}, /* 0xb9f3 */
            {8'h00}, /* 0xb9f2 */
            {8'h00}, /* 0xb9f1 */
            {8'h00}, /* 0xb9f0 */
            {8'h00}, /* 0xb9ef */
            {8'h00}, /* 0xb9ee */
            {8'h00}, /* 0xb9ed */
            {8'h00}, /* 0xb9ec */
            {8'h00}, /* 0xb9eb */
            {8'h00}, /* 0xb9ea */
            {8'h00}, /* 0xb9e9 */
            {8'h00}, /* 0xb9e8 */
            {8'h00}, /* 0xb9e7 */
            {8'h00}, /* 0xb9e6 */
            {8'h00}, /* 0xb9e5 */
            {8'h00}, /* 0xb9e4 */
            {8'h00}, /* 0xb9e3 */
            {8'h00}, /* 0xb9e2 */
            {8'h00}, /* 0xb9e1 */
            {8'h00}, /* 0xb9e0 */
            {8'h00}, /* 0xb9df */
            {8'h00}, /* 0xb9de */
            {8'h00}, /* 0xb9dd */
            {8'h00}, /* 0xb9dc */
            {8'h00}, /* 0xb9db */
            {8'h00}, /* 0xb9da */
            {8'h00}, /* 0xb9d9 */
            {8'h00}, /* 0xb9d8 */
            {8'h00}, /* 0xb9d7 */
            {8'h00}, /* 0xb9d6 */
            {8'h00}, /* 0xb9d5 */
            {8'h00}, /* 0xb9d4 */
            {8'h00}, /* 0xb9d3 */
            {8'h00}, /* 0xb9d2 */
            {8'h00}, /* 0xb9d1 */
            {8'h00}, /* 0xb9d0 */
            {8'h00}, /* 0xb9cf */
            {8'h00}, /* 0xb9ce */
            {8'h00}, /* 0xb9cd */
            {8'h00}, /* 0xb9cc */
            {8'h00}, /* 0xb9cb */
            {8'h00}, /* 0xb9ca */
            {8'h00}, /* 0xb9c9 */
            {8'h00}, /* 0xb9c8 */
            {8'h00}, /* 0xb9c7 */
            {8'h00}, /* 0xb9c6 */
            {8'h00}, /* 0xb9c5 */
            {8'h00}, /* 0xb9c4 */
            {8'h00}, /* 0xb9c3 */
            {8'h00}, /* 0xb9c2 */
            {8'h00}, /* 0xb9c1 */
            {8'h00}, /* 0xb9c0 */
            {8'h00}, /* 0xb9bf */
            {8'h00}, /* 0xb9be */
            {8'h00}, /* 0xb9bd */
            {8'h00}, /* 0xb9bc */
            {8'h00}, /* 0xb9bb */
            {8'h00}, /* 0xb9ba */
            {8'h00}, /* 0xb9b9 */
            {8'h00}, /* 0xb9b8 */
            {8'h00}, /* 0xb9b7 */
            {8'h00}, /* 0xb9b6 */
            {8'h00}, /* 0xb9b5 */
            {8'h00}, /* 0xb9b4 */
            {8'h00}, /* 0xb9b3 */
            {8'h00}, /* 0xb9b2 */
            {8'h00}, /* 0xb9b1 */
            {8'h00}, /* 0xb9b0 */
            {8'h00}, /* 0xb9af */
            {8'h00}, /* 0xb9ae */
            {8'h00}, /* 0xb9ad */
            {8'h00}, /* 0xb9ac */
            {8'h00}, /* 0xb9ab */
            {8'h00}, /* 0xb9aa */
            {8'h00}, /* 0xb9a9 */
            {8'h00}, /* 0xb9a8 */
            {8'h00}, /* 0xb9a7 */
            {8'h00}, /* 0xb9a6 */
            {8'h00}, /* 0xb9a5 */
            {8'h00}, /* 0xb9a4 */
            {8'h00}, /* 0xb9a3 */
            {8'h00}, /* 0xb9a2 */
            {8'h00}, /* 0xb9a1 */
            {8'h00}, /* 0xb9a0 */
            {8'h00}, /* 0xb99f */
            {8'h00}, /* 0xb99e */
            {8'h00}, /* 0xb99d */
            {8'h00}, /* 0xb99c */
            {8'h00}, /* 0xb99b */
            {8'h00}, /* 0xb99a */
            {8'h00}, /* 0xb999 */
            {8'h00}, /* 0xb998 */
            {8'h00}, /* 0xb997 */
            {8'h00}, /* 0xb996 */
            {8'h00}, /* 0xb995 */
            {8'h00}, /* 0xb994 */
            {8'h00}, /* 0xb993 */
            {8'h00}, /* 0xb992 */
            {8'h00}, /* 0xb991 */
            {8'h00}, /* 0xb990 */
            {8'h00}, /* 0xb98f */
            {8'h00}, /* 0xb98e */
            {8'h00}, /* 0xb98d */
            {8'h00}, /* 0xb98c */
            {8'h00}, /* 0xb98b */
            {8'h00}, /* 0xb98a */
            {8'h00}, /* 0xb989 */
            {8'h00}, /* 0xb988 */
            {8'h00}, /* 0xb987 */
            {8'h00}, /* 0xb986 */
            {8'h00}, /* 0xb985 */
            {8'h00}, /* 0xb984 */
            {8'h00}, /* 0xb983 */
            {8'h00}, /* 0xb982 */
            {8'h00}, /* 0xb981 */
            {8'h00}, /* 0xb980 */
            {8'h00}, /* 0xb97f */
            {8'h00}, /* 0xb97e */
            {8'h00}, /* 0xb97d */
            {8'h00}, /* 0xb97c */
            {8'h00}, /* 0xb97b */
            {8'h00}, /* 0xb97a */
            {8'h00}, /* 0xb979 */
            {8'h00}, /* 0xb978 */
            {8'h00}, /* 0xb977 */
            {8'h00}, /* 0xb976 */
            {8'h00}, /* 0xb975 */
            {8'h00}, /* 0xb974 */
            {8'h00}, /* 0xb973 */
            {8'h00}, /* 0xb972 */
            {8'h00}, /* 0xb971 */
            {8'h00}, /* 0xb970 */
            {8'h00}, /* 0xb96f */
            {8'h00}, /* 0xb96e */
            {8'h00}, /* 0xb96d */
            {8'h00}, /* 0xb96c */
            {8'h00}, /* 0xb96b */
            {8'h00}, /* 0xb96a */
            {8'h00}, /* 0xb969 */
            {8'h00}, /* 0xb968 */
            {8'h00}, /* 0xb967 */
            {8'h00}, /* 0xb966 */
            {8'h00}, /* 0xb965 */
            {8'h00}, /* 0xb964 */
            {8'h00}, /* 0xb963 */
            {8'h00}, /* 0xb962 */
            {8'h00}, /* 0xb961 */
            {8'h00}, /* 0xb960 */
            {8'h00}, /* 0xb95f */
            {8'h00}, /* 0xb95e */
            {8'h00}, /* 0xb95d */
            {8'h00}, /* 0xb95c */
            {8'h00}, /* 0xb95b */
            {8'h00}, /* 0xb95a */
            {8'h00}, /* 0xb959 */
            {8'h00}, /* 0xb958 */
            {8'h00}, /* 0xb957 */
            {8'h00}, /* 0xb956 */
            {8'h00}, /* 0xb955 */
            {8'h00}, /* 0xb954 */
            {8'h00}, /* 0xb953 */
            {8'h00}, /* 0xb952 */
            {8'h00}, /* 0xb951 */
            {8'h00}, /* 0xb950 */
            {8'h00}, /* 0xb94f */
            {8'h00}, /* 0xb94e */
            {8'h00}, /* 0xb94d */
            {8'h00}, /* 0xb94c */
            {8'h00}, /* 0xb94b */
            {8'h00}, /* 0xb94a */
            {8'h00}, /* 0xb949 */
            {8'h00}, /* 0xb948 */
            {8'h00}, /* 0xb947 */
            {8'h00}, /* 0xb946 */
            {8'h00}, /* 0xb945 */
            {8'h00}, /* 0xb944 */
            {8'h00}, /* 0xb943 */
            {8'h00}, /* 0xb942 */
            {8'h00}, /* 0xb941 */
            {8'h00}, /* 0xb940 */
            {8'h00}, /* 0xb93f */
            {8'h00}, /* 0xb93e */
            {8'h00}, /* 0xb93d */
            {8'h00}, /* 0xb93c */
            {8'h00}, /* 0xb93b */
            {8'h00}, /* 0xb93a */
            {8'h00}, /* 0xb939 */
            {8'h00}, /* 0xb938 */
            {8'h00}, /* 0xb937 */
            {8'h00}, /* 0xb936 */
            {8'h00}, /* 0xb935 */
            {8'h00}, /* 0xb934 */
            {8'h00}, /* 0xb933 */
            {8'h00}, /* 0xb932 */
            {8'h00}, /* 0xb931 */
            {8'h00}, /* 0xb930 */
            {8'h00}, /* 0xb92f */
            {8'h00}, /* 0xb92e */
            {8'h00}, /* 0xb92d */
            {8'h00}, /* 0xb92c */
            {8'h00}, /* 0xb92b */
            {8'h00}, /* 0xb92a */
            {8'h00}, /* 0xb929 */
            {8'h00}, /* 0xb928 */
            {8'h00}, /* 0xb927 */
            {8'h00}, /* 0xb926 */
            {8'h00}, /* 0xb925 */
            {8'h00}, /* 0xb924 */
            {8'h00}, /* 0xb923 */
            {8'h00}, /* 0xb922 */
            {8'h00}, /* 0xb921 */
            {8'h00}, /* 0xb920 */
            {8'h00}, /* 0xb91f */
            {8'h00}, /* 0xb91e */
            {8'h00}, /* 0xb91d */
            {8'h00}, /* 0xb91c */
            {8'h00}, /* 0xb91b */
            {8'h00}, /* 0xb91a */
            {8'h00}, /* 0xb919 */
            {8'h00}, /* 0xb918 */
            {8'h00}, /* 0xb917 */
            {8'h00}, /* 0xb916 */
            {8'h00}, /* 0xb915 */
            {8'h00}, /* 0xb914 */
            {8'h00}, /* 0xb913 */
            {8'h00}, /* 0xb912 */
            {8'h00}, /* 0xb911 */
            {8'h00}, /* 0xb910 */
            {8'h00}, /* 0xb90f */
            {8'h00}, /* 0xb90e */
            {8'h00}, /* 0xb90d */
            {8'h00}, /* 0xb90c */
            {8'h00}, /* 0xb90b */
            {8'h00}, /* 0xb90a */
            {8'h00}, /* 0xb909 */
            {8'h00}, /* 0xb908 */
            {8'h00}, /* 0xb907 */
            {8'h00}, /* 0xb906 */
            {8'h00}, /* 0xb905 */
            {8'h00}, /* 0xb904 */
            {8'h00}, /* 0xb903 */
            {8'h00}, /* 0xb902 */
            {8'h00}, /* 0xb901 */
            {8'h00}, /* 0xb900 */
            {8'h00}, /* 0xb8ff */
            {8'h00}, /* 0xb8fe */
            {8'h00}, /* 0xb8fd */
            {8'h00}, /* 0xb8fc */
            {8'h00}, /* 0xb8fb */
            {8'h00}, /* 0xb8fa */
            {8'h00}, /* 0xb8f9 */
            {8'h00}, /* 0xb8f8 */
            {8'h00}, /* 0xb8f7 */
            {8'h00}, /* 0xb8f6 */
            {8'h00}, /* 0xb8f5 */
            {8'h00}, /* 0xb8f4 */
            {8'h00}, /* 0xb8f3 */
            {8'h00}, /* 0xb8f2 */
            {8'h00}, /* 0xb8f1 */
            {8'h00}, /* 0xb8f0 */
            {8'h00}, /* 0xb8ef */
            {8'h00}, /* 0xb8ee */
            {8'h00}, /* 0xb8ed */
            {8'h00}, /* 0xb8ec */
            {8'h00}, /* 0xb8eb */
            {8'h00}, /* 0xb8ea */
            {8'h00}, /* 0xb8e9 */
            {8'h00}, /* 0xb8e8 */
            {8'h00}, /* 0xb8e7 */
            {8'h00}, /* 0xb8e6 */
            {8'h00}, /* 0xb8e5 */
            {8'h00}, /* 0xb8e4 */
            {8'h00}, /* 0xb8e3 */
            {8'h00}, /* 0xb8e2 */
            {8'h00}, /* 0xb8e1 */
            {8'h00}, /* 0xb8e0 */
            {8'h00}, /* 0xb8df */
            {8'h00}, /* 0xb8de */
            {8'h00}, /* 0xb8dd */
            {8'h00}, /* 0xb8dc */
            {8'h00}, /* 0xb8db */
            {8'h00}, /* 0xb8da */
            {8'h00}, /* 0xb8d9 */
            {8'h00}, /* 0xb8d8 */
            {8'h00}, /* 0xb8d7 */
            {8'h00}, /* 0xb8d6 */
            {8'h00}, /* 0xb8d5 */
            {8'h00}, /* 0xb8d4 */
            {8'h00}, /* 0xb8d3 */
            {8'h00}, /* 0xb8d2 */
            {8'h00}, /* 0xb8d1 */
            {8'h00}, /* 0xb8d0 */
            {8'h00}, /* 0xb8cf */
            {8'h00}, /* 0xb8ce */
            {8'h00}, /* 0xb8cd */
            {8'h00}, /* 0xb8cc */
            {8'h00}, /* 0xb8cb */
            {8'h00}, /* 0xb8ca */
            {8'h00}, /* 0xb8c9 */
            {8'h00}, /* 0xb8c8 */
            {8'h00}, /* 0xb8c7 */
            {8'h00}, /* 0xb8c6 */
            {8'h00}, /* 0xb8c5 */
            {8'h00}, /* 0xb8c4 */
            {8'h00}, /* 0xb8c3 */
            {8'h00}, /* 0xb8c2 */
            {8'h00}, /* 0xb8c1 */
            {8'h00}, /* 0xb8c0 */
            {8'h00}, /* 0xb8bf */
            {8'h00}, /* 0xb8be */
            {8'h00}, /* 0xb8bd */
            {8'h00}, /* 0xb8bc */
            {8'h00}, /* 0xb8bb */
            {8'h00}, /* 0xb8ba */
            {8'h00}, /* 0xb8b9 */
            {8'h00}, /* 0xb8b8 */
            {8'h00}, /* 0xb8b7 */
            {8'h00}, /* 0xb8b6 */
            {8'h00}, /* 0xb8b5 */
            {8'h00}, /* 0xb8b4 */
            {8'h00}, /* 0xb8b3 */
            {8'h00}, /* 0xb8b2 */
            {8'h00}, /* 0xb8b1 */
            {8'h00}, /* 0xb8b0 */
            {8'h00}, /* 0xb8af */
            {8'h00}, /* 0xb8ae */
            {8'h00}, /* 0xb8ad */
            {8'h00}, /* 0xb8ac */
            {8'h00}, /* 0xb8ab */
            {8'h00}, /* 0xb8aa */
            {8'h00}, /* 0xb8a9 */
            {8'h00}, /* 0xb8a8 */
            {8'h00}, /* 0xb8a7 */
            {8'h00}, /* 0xb8a6 */
            {8'h00}, /* 0xb8a5 */
            {8'h00}, /* 0xb8a4 */
            {8'h00}, /* 0xb8a3 */
            {8'h00}, /* 0xb8a2 */
            {8'h00}, /* 0xb8a1 */
            {8'h00}, /* 0xb8a0 */
            {8'h00}, /* 0xb89f */
            {8'h00}, /* 0xb89e */
            {8'h00}, /* 0xb89d */
            {8'h00}, /* 0xb89c */
            {8'h00}, /* 0xb89b */
            {8'h00}, /* 0xb89a */
            {8'h00}, /* 0xb899 */
            {8'h00}, /* 0xb898 */
            {8'h00}, /* 0xb897 */
            {8'h00}, /* 0xb896 */
            {8'h00}, /* 0xb895 */
            {8'h00}, /* 0xb894 */
            {8'h00}, /* 0xb893 */
            {8'h00}, /* 0xb892 */
            {8'h00}, /* 0xb891 */
            {8'h00}, /* 0xb890 */
            {8'h00}, /* 0xb88f */
            {8'h00}, /* 0xb88e */
            {8'h00}, /* 0xb88d */
            {8'h00}, /* 0xb88c */
            {8'h00}, /* 0xb88b */
            {8'h00}, /* 0xb88a */
            {8'h00}, /* 0xb889 */
            {8'h00}, /* 0xb888 */
            {8'h00}, /* 0xb887 */
            {8'h00}, /* 0xb886 */
            {8'h00}, /* 0xb885 */
            {8'h00}, /* 0xb884 */
            {8'h00}, /* 0xb883 */
            {8'h00}, /* 0xb882 */
            {8'h00}, /* 0xb881 */
            {8'h00}, /* 0xb880 */
            {8'h00}, /* 0xb87f */
            {8'h00}, /* 0xb87e */
            {8'h00}, /* 0xb87d */
            {8'h00}, /* 0xb87c */
            {8'h00}, /* 0xb87b */
            {8'h00}, /* 0xb87a */
            {8'h00}, /* 0xb879 */
            {8'h00}, /* 0xb878 */
            {8'h00}, /* 0xb877 */
            {8'h00}, /* 0xb876 */
            {8'h00}, /* 0xb875 */
            {8'h00}, /* 0xb874 */
            {8'h00}, /* 0xb873 */
            {8'h00}, /* 0xb872 */
            {8'h00}, /* 0xb871 */
            {8'h00}, /* 0xb870 */
            {8'h00}, /* 0xb86f */
            {8'h00}, /* 0xb86e */
            {8'h00}, /* 0xb86d */
            {8'h00}, /* 0xb86c */
            {8'h00}, /* 0xb86b */
            {8'h00}, /* 0xb86a */
            {8'h00}, /* 0xb869 */
            {8'h00}, /* 0xb868 */
            {8'h00}, /* 0xb867 */
            {8'h00}, /* 0xb866 */
            {8'h00}, /* 0xb865 */
            {8'h00}, /* 0xb864 */
            {8'h00}, /* 0xb863 */
            {8'h00}, /* 0xb862 */
            {8'h00}, /* 0xb861 */
            {8'h00}, /* 0xb860 */
            {8'h00}, /* 0xb85f */
            {8'h00}, /* 0xb85e */
            {8'h00}, /* 0xb85d */
            {8'h00}, /* 0xb85c */
            {8'h00}, /* 0xb85b */
            {8'h00}, /* 0xb85a */
            {8'h00}, /* 0xb859 */
            {8'h00}, /* 0xb858 */
            {8'h00}, /* 0xb857 */
            {8'h00}, /* 0xb856 */
            {8'h00}, /* 0xb855 */
            {8'h00}, /* 0xb854 */
            {8'h00}, /* 0xb853 */
            {8'h00}, /* 0xb852 */
            {8'h00}, /* 0xb851 */
            {8'h00}, /* 0xb850 */
            {8'h00}, /* 0xb84f */
            {8'h00}, /* 0xb84e */
            {8'h00}, /* 0xb84d */
            {8'h00}, /* 0xb84c */
            {8'h00}, /* 0xb84b */
            {8'h00}, /* 0xb84a */
            {8'h00}, /* 0xb849 */
            {8'h00}, /* 0xb848 */
            {8'h00}, /* 0xb847 */
            {8'h00}, /* 0xb846 */
            {8'h00}, /* 0xb845 */
            {8'h00}, /* 0xb844 */
            {8'h00}, /* 0xb843 */
            {8'h00}, /* 0xb842 */
            {8'h00}, /* 0xb841 */
            {8'h00}, /* 0xb840 */
            {8'h00}, /* 0xb83f */
            {8'h00}, /* 0xb83e */
            {8'h00}, /* 0xb83d */
            {8'h00}, /* 0xb83c */
            {8'h00}, /* 0xb83b */
            {8'h00}, /* 0xb83a */
            {8'h00}, /* 0xb839 */
            {8'h00}, /* 0xb838 */
            {8'h00}, /* 0xb837 */
            {8'h00}, /* 0xb836 */
            {8'h00}, /* 0xb835 */
            {8'h00}, /* 0xb834 */
            {8'h00}, /* 0xb833 */
            {8'h00}, /* 0xb832 */
            {8'h00}, /* 0xb831 */
            {8'h00}, /* 0xb830 */
            {8'h00}, /* 0xb82f */
            {8'h00}, /* 0xb82e */
            {8'h00}, /* 0xb82d */
            {8'h00}, /* 0xb82c */
            {8'h00}, /* 0xb82b */
            {8'h00}, /* 0xb82a */
            {8'h00}, /* 0xb829 */
            {8'h00}, /* 0xb828 */
            {8'h00}, /* 0xb827 */
            {8'h00}, /* 0xb826 */
            {8'h00}, /* 0xb825 */
            {8'h00}, /* 0xb824 */
            {8'h00}, /* 0xb823 */
            {8'h00}, /* 0xb822 */
            {8'h00}, /* 0xb821 */
            {8'h00}, /* 0xb820 */
            {8'h00}, /* 0xb81f */
            {8'h00}, /* 0xb81e */
            {8'h00}, /* 0xb81d */
            {8'h00}, /* 0xb81c */
            {8'h00}, /* 0xb81b */
            {8'h00}, /* 0xb81a */
            {8'h00}, /* 0xb819 */
            {8'h00}, /* 0xb818 */
            {8'h00}, /* 0xb817 */
            {8'h00}, /* 0xb816 */
            {8'h00}, /* 0xb815 */
            {8'h00}, /* 0xb814 */
            {8'h00}, /* 0xb813 */
            {8'h00}, /* 0xb812 */
            {8'h00}, /* 0xb811 */
            {8'h00}, /* 0xb810 */
            {8'h00}, /* 0xb80f */
            {8'h00}, /* 0xb80e */
            {8'h00}, /* 0xb80d */
            {8'h00}, /* 0xb80c */
            {8'h00}, /* 0xb80b */
            {8'h00}, /* 0xb80a */
            {8'h00}, /* 0xb809 */
            {8'h00}, /* 0xb808 */
            {8'h00}, /* 0xb807 */
            {8'h00}, /* 0xb806 */
            {8'h00}, /* 0xb805 */
            {8'h00}, /* 0xb804 */
            {8'h00}, /* 0xb803 */
            {8'h00}, /* 0xb802 */
            {8'h00}, /* 0xb801 */
            {8'h00}, /* 0xb800 */
            {8'h00}, /* 0xb7ff */
            {8'h00}, /* 0xb7fe */
            {8'h00}, /* 0xb7fd */
            {8'h00}, /* 0xb7fc */
            {8'h00}, /* 0xb7fb */
            {8'h00}, /* 0xb7fa */
            {8'h00}, /* 0xb7f9 */
            {8'h00}, /* 0xb7f8 */
            {8'h00}, /* 0xb7f7 */
            {8'h00}, /* 0xb7f6 */
            {8'h00}, /* 0xb7f5 */
            {8'h00}, /* 0xb7f4 */
            {8'h00}, /* 0xb7f3 */
            {8'h00}, /* 0xb7f2 */
            {8'h00}, /* 0xb7f1 */
            {8'h00}, /* 0xb7f0 */
            {8'h00}, /* 0xb7ef */
            {8'h00}, /* 0xb7ee */
            {8'h00}, /* 0xb7ed */
            {8'h00}, /* 0xb7ec */
            {8'h00}, /* 0xb7eb */
            {8'h00}, /* 0xb7ea */
            {8'h00}, /* 0xb7e9 */
            {8'h00}, /* 0xb7e8 */
            {8'h00}, /* 0xb7e7 */
            {8'h00}, /* 0xb7e6 */
            {8'h00}, /* 0xb7e5 */
            {8'h00}, /* 0xb7e4 */
            {8'h00}, /* 0xb7e3 */
            {8'h00}, /* 0xb7e2 */
            {8'h00}, /* 0xb7e1 */
            {8'h00}, /* 0xb7e0 */
            {8'h00}, /* 0xb7df */
            {8'h00}, /* 0xb7de */
            {8'h00}, /* 0xb7dd */
            {8'h00}, /* 0xb7dc */
            {8'h00}, /* 0xb7db */
            {8'h00}, /* 0xb7da */
            {8'h00}, /* 0xb7d9 */
            {8'h00}, /* 0xb7d8 */
            {8'h00}, /* 0xb7d7 */
            {8'h00}, /* 0xb7d6 */
            {8'h00}, /* 0xb7d5 */
            {8'h00}, /* 0xb7d4 */
            {8'h00}, /* 0xb7d3 */
            {8'h00}, /* 0xb7d2 */
            {8'h00}, /* 0xb7d1 */
            {8'h00}, /* 0xb7d0 */
            {8'h00}, /* 0xb7cf */
            {8'h00}, /* 0xb7ce */
            {8'h00}, /* 0xb7cd */
            {8'h00}, /* 0xb7cc */
            {8'h00}, /* 0xb7cb */
            {8'h00}, /* 0xb7ca */
            {8'h00}, /* 0xb7c9 */
            {8'h00}, /* 0xb7c8 */
            {8'h00}, /* 0xb7c7 */
            {8'h00}, /* 0xb7c6 */
            {8'h00}, /* 0xb7c5 */
            {8'h00}, /* 0xb7c4 */
            {8'h00}, /* 0xb7c3 */
            {8'h00}, /* 0xb7c2 */
            {8'h00}, /* 0xb7c1 */
            {8'h00}, /* 0xb7c0 */
            {8'h00}, /* 0xb7bf */
            {8'h00}, /* 0xb7be */
            {8'h00}, /* 0xb7bd */
            {8'h00}, /* 0xb7bc */
            {8'h00}, /* 0xb7bb */
            {8'h00}, /* 0xb7ba */
            {8'h00}, /* 0xb7b9 */
            {8'h00}, /* 0xb7b8 */
            {8'h00}, /* 0xb7b7 */
            {8'h00}, /* 0xb7b6 */
            {8'h00}, /* 0xb7b5 */
            {8'h00}, /* 0xb7b4 */
            {8'h00}, /* 0xb7b3 */
            {8'h00}, /* 0xb7b2 */
            {8'h00}, /* 0xb7b1 */
            {8'h00}, /* 0xb7b0 */
            {8'h00}, /* 0xb7af */
            {8'h00}, /* 0xb7ae */
            {8'h00}, /* 0xb7ad */
            {8'h00}, /* 0xb7ac */
            {8'h00}, /* 0xb7ab */
            {8'h00}, /* 0xb7aa */
            {8'h00}, /* 0xb7a9 */
            {8'h00}, /* 0xb7a8 */
            {8'h00}, /* 0xb7a7 */
            {8'h00}, /* 0xb7a6 */
            {8'h00}, /* 0xb7a5 */
            {8'h00}, /* 0xb7a4 */
            {8'h00}, /* 0xb7a3 */
            {8'h00}, /* 0xb7a2 */
            {8'h00}, /* 0xb7a1 */
            {8'h00}, /* 0xb7a0 */
            {8'h00}, /* 0xb79f */
            {8'h00}, /* 0xb79e */
            {8'h00}, /* 0xb79d */
            {8'h00}, /* 0xb79c */
            {8'h00}, /* 0xb79b */
            {8'h00}, /* 0xb79a */
            {8'h00}, /* 0xb799 */
            {8'h00}, /* 0xb798 */
            {8'h00}, /* 0xb797 */
            {8'h00}, /* 0xb796 */
            {8'h00}, /* 0xb795 */
            {8'h00}, /* 0xb794 */
            {8'h00}, /* 0xb793 */
            {8'h00}, /* 0xb792 */
            {8'h00}, /* 0xb791 */
            {8'h00}, /* 0xb790 */
            {8'h00}, /* 0xb78f */
            {8'h00}, /* 0xb78e */
            {8'h00}, /* 0xb78d */
            {8'h00}, /* 0xb78c */
            {8'h00}, /* 0xb78b */
            {8'h00}, /* 0xb78a */
            {8'h00}, /* 0xb789 */
            {8'h00}, /* 0xb788 */
            {8'h00}, /* 0xb787 */
            {8'h00}, /* 0xb786 */
            {8'h00}, /* 0xb785 */
            {8'h00}, /* 0xb784 */
            {8'h00}, /* 0xb783 */
            {8'h00}, /* 0xb782 */
            {8'h00}, /* 0xb781 */
            {8'h00}, /* 0xb780 */
            {8'h00}, /* 0xb77f */
            {8'h00}, /* 0xb77e */
            {8'h00}, /* 0xb77d */
            {8'h00}, /* 0xb77c */
            {8'h00}, /* 0xb77b */
            {8'h00}, /* 0xb77a */
            {8'h00}, /* 0xb779 */
            {8'h00}, /* 0xb778 */
            {8'h00}, /* 0xb777 */
            {8'h00}, /* 0xb776 */
            {8'h00}, /* 0xb775 */
            {8'h00}, /* 0xb774 */
            {8'h00}, /* 0xb773 */
            {8'h00}, /* 0xb772 */
            {8'h00}, /* 0xb771 */
            {8'h00}, /* 0xb770 */
            {8'h00}, /* 0xb76f */
            {8'h00}, /* 0xb76e */
            {8'h00}, /* 0xb76d */
            {8'h00}, /* 0xb76c */
            {8'h00}, /* 0xb76b */
            {8'h00}, /* 0xb76a */
            {8'h00}, /* 0xb769 */
            {8'h00}, /* 0xb768 */
            {8'h00}, /* 0xb767 */
            {8'h00}, /* 0xb766 */
            {8'h00}, /* 0xb765 */
            {8'h00}, /* 0xb764 */
            {8'h00}, /* 0xb763 */
            {8'h00}, /* 0xb762 */
            {8'h00}, /* 0xb761 */
            {8'h00}, /* 0xb760 */
            {8'h00}, /* 0xb75f */
            {8'h00}, /* 0xb75e */
            {8'h00}, /* 0xb75d */
            {8'h00}, /* 0xb75c */
            {8'h00}, /* 0xb75b */
            {8'h00}, /* 0xb75a */
            {8'h00}, /* 0xb759 */
            {8'h00}, /* 0xb758 */
            {8'h00}, /* 0xb757 */
            {8'h00}, /* 0xb756 */
            {8'h00}, /* 0xb755 */
            {8'h00}, /* 0xb754 */
            {8'h00}, /* 0xb753 */
            {8'h00}, /* 0xb752 */
            {8'h00}, /* 0xb751 */
            {8'h00}, /* 0xb750 */
            {8'h00}, /* 0xb74f */
            {8'h00}, /* 0xb74e */
            {8'h00}, /* 0xb74d */
            {8'h00}, /* 0xb74c */
            {8'h00}, /* 0xb74b */
            {8'h00}, /* 0xb74a */
            {8'h00}, /* 0xb749 */
            {8'h00}, /* 0xb748 */
            {8'h00}, /* 0xb747 */
            {8'h00}, /* 0xb746 */
            {8'h00}, /* 0xb745 */
            {8'h00}, /* 0xb744 */
            {8'h00}, /* 0xb743 */
            {8'h00}, /* 0xb742 */
            {8'h00}, /* 0xb741 */
            {8'h00}, /* 0xb740 */
            {8'h00}, /* 0xb73f */
            {8'h00}, /* 0xb73e */
            {8'h00}, /* 0xb73d */
            {8'h00}, /* 0xb73c */
            {8'h00}, /* 0xb73b */
            {8'h00}, /* 0xb73a */
            {8'h00}, /* 0xb739 */
            {8'h00}, /* 0xb738 */
            {8'h00}, /* 0xb737 */
            {8'h00}, /* 0xb736 */
            {8'h00}, /* 0xb735 */
            {8'h00}, /* 0xb734 */
            {8'h00}, /* 0xb733 */
            {8'h00}, /* 0xb732 */
            {8'h00}, /* 0xb731 */
            {8'h00}, /* 0xb730 */
            {8'h00}, /* 0xb72f */
            {8'h00}, /* 0xb72e */
            {8'h00}, /* 0xb72d */
            {8'h00}, /* 0xb72c */
            {8'h00}, /* 0xb72b */
            {8'h00}, /* 0xb72a */
            {8'h00}, /* 0xb729 */
            {8'h00}, /* 0xb728 */
            {8'h00}, /* 0xb727 */
            {8'h00}, /* 0xb726 */
            {8'h00}, /* 0xb725 */
            {8'h00}, /* 0xb724 */
            {8'h00}, /* 0xb723 */
            {8'h00}, /* 0xb722 */
            {8'h00}, /* 0xb721 */
            {8'h00}, /* 0xb720 */
            {8'h00}, /* 0xb71f */
            {8'h00}, /* 0xb71e */
            {8'h00}, /* 0xb71d */
            {8'h00}, /* 0xb71c */
            {8'h00}, /* 0xb71b */
            {8'h00}, /* 0xb71a */
            {8'h00}, /* 0xb719 */
            {8'h00}, /* 0xb718 */
            {8'h00}, /* 0xb717 */
            {8'h00}, /* 0xb716 */
            {8'h00}, /* 0xb715 */
            {8'h00}, /* 0xb714 */
            {8'h00}, /* 0xb713 */
            {8'h00}, /* 0xb712 */
            {8'h00}, /* 0xb711 */
            {8'h00}, /* 0xb710 */
            {8'h00}, /* 0xb70f */
            {8'h00}, /* 0xb70e */
            {8'h00}, /* 0xb70d */
            {8'h00}, /* 0xb70c */
            {8'h00}, /* 0xb70b */
            {8'h00}, /* 0xb70a */
            {8'h00}, /* 0xb709 */
            {8'h00}, /* 0xb708 */
            {8'h00}, /* 0xb707 */
            {8'h00}, /* 0xb706 */
            {8'h00}, /* 0xb705 */
            {8'h00}, /* 0xb704 */
            {8'h00}, /* 0xb703 */
            {8'h00}, /* 0xb702 */
            {8'h00}, /* 0xb701 */
            {8'h00}, /* 0xb700 */
            {8'h00}, /* 0xb6ff */
            {8'h00}, /* 0xb6fe */
            {8'h00}, /* 0xb6fd */
            {8'h00}, /* 0xb6fc */
            {8'h00}, /* 0xb6fb */
            {8'h00}, /* 0xb6fa */
            {8'h00}, /* 0xb6f9 */
            {8'h00}, /* 0xb6f8 */
            {8'h00}, /* 0xb6f7 */
            {8'h00}, /* 0xb6f6 */
            {8'h00}, /* 0xb6f5 */
            {8'h00}, /* 0xb6f4 */
            {8'h00}, /* 0xb6f3 */
            {8'h00}, /* 0xb6f2 */
            {8'h00}, /* 0xb6f1 */
            {8'h00}, /* 0xb6f0 */
            {8'h00}, /* 0xb6ef */
            {8'h00}, /* 0xb6ee */
            {8'h00}, /* 0xb6ed */
            {8'h00}, /* 0xb6ec */
            {8'h00}, /* 0xb6eb */
            {8'h00}, /* 0xb6ea */
            {8'h00}, /* 0xb6e9 */
            {8'h00}, /* 0xb6e8 */
            {8'h00}, /* 0xb6e7 */
            {8'h00}, /* 0xb6e6 */
            {8'h00}, /* 0xb6e5 */
            {8'h00}, /* 0xb6e4 */
            {8'h00}, /* 0xb6e3 */
            {8'h00}, /* 0xb6e2 */
            {8'h00}, /* 0xb6e1 */
            {8'h00}, /* 0xb6e0 */
            {8'h00}, /* 0xb6df */
            {8'h00}, /* 0xb6de */
            {8'h00}, /* 0xb6dd */
            {8'h00}, /* 0xb6dc */
            {8'h00}, /* 0xb6db */
            {8'h00}, /* 0xb6da */
            {8'h00}, /* 0xb6d9 */
            {8'h00}, /* 0xb6d8 */
            {8'h00}, /* 0xb6d7 */
            {8'h00}, /* 0xb6d6 */
            {8'h00}, /* 0xb6d5 */
            {8'h00}, /* 0xb6d4 */
            {8'h00}, /* 0xb6d3 */
            {8'h00}, /* 0xb6d2 */
            {8'h00}, /* 0xb6d1 */
            {8'h00}, /* 0xb6d0 */
            {8'h00}, /* 0xb6cf */
            {8'h00}, /* 0xb6ce */
            {8'h00}, /* 0xb6cd */
            {8'h00}, /* 0xb6cc */
            {8'h00}, /* 0xb6cb */
            {8'h00}, /* 0xb6ca */
            {8'h00}, /* 0xb6c9 */
            {8'h00}, /* 0xb6c8 */
            {8'h00}, /* 0xb6c7 */
            {8'h00}, /* 0xb6c6 */
            {8'h00}, /* 0xb6c5 */
            {8'h00}, /* 0xb6c4 */
            {8'h00}, /* 0xb6c3 */
            {8'h00}, /* 0xb6c2 */
            {8'h00}, /* 0xb6c1 */
            {8'h00}, /* 0xb6c0 */
            {8'h00}, /* 0xb6bf */
            {8'h00}, /* 0xb6be */
            {8'h00}, /* 0xb6bd */
            {8'h00}, /* 0xb6bc */
            {8'h00}, /* 0xb6bb */
            {8'h00}, /* 0xb6ba */
            {8'h00}, /* 0xb6b9 */
            {8'h00}, /* 0xb6b8 */
            {8'h00}, /* 0xb6b7 */
            {8'h00}, /* 0xb6b6 */
            {8'h00}, /* 0xb6b5 */
            {8'h00}, /* 0xb6b4 */
            {8'h00}, /* 0xb6b3 */
            {8'h00}, /* 0xb6b2 */
            {8'h00}, /* 0xb6b1 */
            {8'h00}, /* 0xb6b0 */
            {8'h00}, /* 0xb6af */
            {8'h00}, /* 0xb6ae */
            {8'h00}, /* 0xb6ad */
            {8'h00}, /* 0xb6ac */
            {8'h00}, /* 0xb6ab */
            {8'h00}, /* 0xb6aa */
            {8'h00}, /* 0xb6a9 */
            {8'h00}, /* 0xb6a8 */
            {8'h00}, /* 0xb6a7 */
            {8'h00}, /* 0xb6a6 */
            {8'h00}, /* 0xb6a5 */
            {8'h00}, /* 0xb6a4 */
            {8'h00}, /* 0xb6a3 */
            {8'h00}, /* 0xb6a2 */
            {8'h00}, /* 0xb6a1 */
            {8'h00}, /* 0xb6a0 */
            {8'h00}, /* 0xb69f */
            {8'h00}, /* 0xb69e */
            {8'h00}, /* 0xb69d */
            {8'h00}, /* 0xb69c */
            {8'h00}, /* 0xb69b */
            {8'h00}, /* 0xb69a */
            {8'h00}, /* 0xb699 */
            {8'h00}, /* 0xb698 */
            {8'h00}, /* 0xb697 */
            {8'h00}, /* 0xb696 */
            {8'h00}, /* 0xb695 */
            {8'h00}, /* 0xb694 */
            {8'h00}, /* 0xb693 */
            {8'h00}, /* 0xb692 */
            {8'h00}, /* 0xb691 */
            {8'h00}, /* 0xb690 */
            {8'h00}, /* 0xb68f */
            {8'h00}, /* 0xb68e */
            {8'h00}, /* 0xb68d */
            {8'h00}, /* 0xb68c */
            {8'h00}, /* 0xb68b */
            {8'h00}, /* 0xb68a */
            {8'h00}, /* 0xb689 */
            {8'h00}, /* 0xb688 */
            {8'h00}, /* 0xb687 */
            {8'h00}, /* 0xb686 */
            {8'h00}, /* 0xb685 */
            {8'h00}, /* 0xb684 */
            {8'h00}, /* 0xb683 */
            {8'h00}, /* 0xb682 */
            {8'h00}, /* 0xb681 */
            {8'h00}, /* 0xb680 */
            {8'h00}, /* 0xb67f */
            {8'h00}, /* 0xb67e */
            {8'h00}, /* 0xb67d */
            {8'h00}, /* 0xb67c */
            {8'h00}, /* 0xb67b */
            {8'h00}, /* 0xb67a */
            {8'h00}, /* 0xb679 */
            {8'h00}, /* 0xb678 */
            {8'h00}, /* 0xb677 */
            {8'h00}, /* 0xb676 */
            {8'h00}, /* 0xb675 */
            {8'h00}, /* 0xb674 */
            {8'h00}, /* 0xb673 */
            {8'h00}, /* 0xb672 */
            {8'h00}, /* 0xb671 */
            {8'h00}, /* 0xb670 */
            {8'h00}, /* 0xb66f */
            {8'h00}, /* 0xb66e */
            {8'h00}, /* 0xb66d */
            {8'h00}, /* 0xb66c */
            {8'h00}, /* 0xb66b */
            {8'h00}, /* 0xb66a */
            {8'h00}, /* 0xb669 */
            {8'h00}, /* 0xb668 */
            {8'h00}, /* 0xb667 */
            {8'h00}, /* 0xb666 */
            {8'h00}, /* 0xb665 */
            {8'h00}, /* 0xb664 */
            {8'h00}, /* 0xb663 */
            {8'h00}, /* 0xb662 */
            {8'h00}, /* 0xb661 */
            {8'h00}, /* 0xb660 */
            {8'h00}, /* 0xb65f */
            {8'h00}, /* 0xb65e */
            {8'h00}, /* 0xb65d */
            {8'h00}, /* 0xb65c */
            {8'h00}, /* 0xb65b */
            {8'h00}, /* 0xb65a */
            {8'h00}, /* 0xb659 */
            {8'h00}, /* 0xb658 */
            {8'h00}, /* 0xb657 */
            {8'h00}, /* 0xb656 */
            {8'h00}, /* 0xb655 */
            {8'h00}, /* 0xb654 */
            {8'h00}, /* 0xb653 */
            {8'h00}, /* 0xb652 */
            {8'h00}, /* 0xb651 */
            {8'h00}, /* 0xb650 */
            {8'h00}, /* 0xb64f */
            {8'h00}, /* 0xb64e */
            {8'h00}, /* 0xb64d */
            {8'h00}, /* 0xb64c */
            {8'h00}, /* 0xb64b */
            {8'h00}, /* 0xb64a */
            {8'h00}, /* 0xb649 */
            {8'h00}, /* 0xb648 */
            {8'h00}, /* 0xb647 */
            {8'h00}, /* 0xb646 */
            {8'h00}, /* 0xb645 */
            {8'h00}, /* 0xb644 */
            {8'h00}, /* 0xb643 */
            {8'h00}, /* 0xb642 */
            {8'h00}, /* 0xb641 */
            {8'h00}, /* 0xb640 */
            {8'h00}, /* 0xb63f */
            {8'h00}, /* 0xb63e */
            {8'h00}, /* 0xb63d */
            {8'h00}, /* 0xb63c */
            {8'h00}, /* 0xb63b */
            {8'h00}, /* 0xb63a */
            {8'h00}, /* 0xb639 */
            {8'h00}, /* 0xb638 */
            {8'h00}, /* 0xb637 */
            {8'h00}, /* 0xb636 */
            {8'h00}, /* 0xb635 */
            {8'h00}, /* 0xb634 */
            {8'h00}, /* 0xb633 */
            {8'h00}, /* 0xb632 */
            {8'h00}, /* 0xb631 */
            {8'h00}, /* 0xb630 */
            {8'h00}, /* 0xb62f */
            {8'h00}, /* 0xb62e */
            {8'h00}, /* 0xb62d */
            {8'h00}, /* 0xb62c */
            {8'h00}, /* 0xb62b */
            {8'h00}, /* 0xb62a */
            {8'h00}, /* 0xb629 */
            {8'h00}, /* 0xb628 */
            {8'h00}, /* 0xb627 */
            {8'h00}, /* 0xb626 */
            {8'h00}, /* 0xb625 */
            {8'h00}, /* 0xb624 */
            {8'h00}, /* 0xb623 */
            {8'h00}, /* 0xb622 */
            {8'h00}, /* 0xb621 */
            {8'h00}, /* 0xb620 */
            {8'h00}, /* 0xb61f */
            {8'h00}, /* 0xb61e */
            {8'h00}, /* 0xb61d */
            {8'h00}, /* 0xb61c */
            {8'h00}, /* 0xb61b */
            {8'h00}, /* 0xb61a */
            {8'h00}, /* 0xb619 */
            {8'h00}, /* 0xb618 */
            {8'h00}, /* 0xb617 */
            {8'h00}, /* 0xb616 */
            {8'h00}, /* 0xb615 */
            {8'h00}, /* 0xb614 */
            {8'h00}, /* 0xb613 */
            {8'h00}, /* 0xb612 */
            {8'h00}, /* 0xb611 */
            {8'h00}, /* 0xb610 */
            {8'h00}, /* 0xb60f */
            {8'h00}, /* 0xb60e */
            {8'h00}, /* 0xb60d */
            {8'h00}, /* 0xb60c */
            {8'h00}, /* 0xb60b */
            {8'h00}, /* 0xb60a */
            {8'h00}, /* 0xb609 */
            {8'h00}, /* 0xb608 */
            {8'h00}, /* 0xb607 */
            {8'h00}, /* 0xb606 */
            {8'h00}, /* 0xb605 */
            {8'h00}, /* 0xb604 */
            {8'h00}, /* 0xb603 */
            {8'h00}, /* 0xb602 */
            {8'h00}, /* 0xb601 */
            {8'h00}, /* 0xb600 */
            {8'h00}, /* 0xb5ff */
            {8'h00}, /* 0xb5fe */
            {8'h00}, /* 0xb5fd */
            {8'h00}, /* 0xb5fc */
            {8'h00}, /* 0xb5fb */
            {8'h00}, /* 0xb5fa */
            {8'h00}, /* 0xb5f9 */
            {8'h00}, /* 0xb5f8 */
            {8'h00}, /* 0xb5f7 */
            {8'h00}, /* 0xb5f6 */
            {8'h00}, /* 0xb5f5 */
            {8'h00}, /* 0xb5f4 */
            {8'h00}, /* 0xb5f3 */
            {8'h00}, /* 0xb5f2 */
            {8'h00}, /* 0xb5f1 */
            {8'h00}, /* 0xb5f0 */
            {8'h00}, /* 0xb5ef */
            {8'h00}, /* 0xb5ee */
            {8'h00}, /* 0xb5ed */
            {8'h00}, /* 0xb5ec */
            {8'h00}, /* 0xb5eb */
            {8'h00}, /* 0xb5ea */
            {8'h00}, /* 0xb5e9 */
            {8'h00}, /* 0xb5e8 */
            {8'h00}, /* 0xb5e7 */
            {8'h00}, /* 0xb5e6 */
            {8'h00}, /* 0xb5e5 */
            {8'h00}, /* 0xb5e4 */
            {8'h00}, /* 0xb5e3 */
            {8'h00}, /* 0xb5e2 */
            {8'h00}, /* 0xb5e1 */
            {8'h00}, /* 0xb5e0 */
            {8'h00}, /* 0xb5df */
            {8'h00}, /* 0xb5de */
            {8'h00}, /* 0xb5dd */
            {8'h00}, /* 0xb5dc */
            {8'h00}, /* 0xb5db */
            {8'h00}, /* 0xb5da */
            {8'h00}, /* 0xb5d9 */
            {8'h00}, /* 0xb5d8 */
            {8'h00}, /* 0xb5d7 */
            {8'h00}, /* 0xb5d6 */
            {8'h00}, /* 0xb5d5 */
            {8'h00}, /* 0xb5d4 */
            {8'h00}, /* 0xb5d3 */
            {8'h00}, /* 0xb5d2 */
            {8'h00}, /* 0xb5d1 */
            {8'h00}, /* 0xb5d0 */
            {8'h00}, /* 0xb5cf */
            {8'h00}, /* 0xb5ce */
            {8'h00}, /* 0xb5cd */
            {8'h00}, /* 0xb5cc */
            {8'h00}, /* 0xb5cb */
            {8'h00}, /* 0xb5ca */
            {8'h00}, /* 0xb5c9 */
            {8'h00}, /* 0xb5c8 */
            {8'h00}, /* 0xb5c7 */
            {8'h00}, /* 0xb5c6 */
            {8'h00}, /* 0xb5c5 */
            {8'h00}, /* 0xb5c4 */
            {8'h00}, /* 0xb5c3 */
            {8'h00}, /* 0xb5c2 */
            {8'h00}, /* 0xb5c1 */
            {8'h00}, /* 0xb5c0 */
            {8'h00}, /* 0xb5bf */
            {8'h00}, /* 0xb5be */
            {8'h00}, /* 0xb5bd */
            {8'h00}, /* 0xb5bc */
            {8'h00}, /* 0xb5bb */
            {8'h00}, /* 0xb5ba */
            {8'h00}, /* 0xb5b9 */
            {8'h00}, /* 0xb5b8 */
            {8'h00}, /* 0xb5b7 */
            {8'h00}, /* 0xb5b6 */
            {8'h00}, /* 0xb5b5 */
            {8'h00}, /* 0xb5b4 */
            {8'h00}, /* 0xb5b3 */
            {8'h00}, /* 0xb5b2 */
            {8'h00}, /* 0xb5b1 */
            {8'h00}, /* 0xb5b0 */
            {8'h00}, /* 0xb5af */
            {8'h00}, /* 0xb5ae */
            {8'h00}, /* 0xb5ad */
            {8'h00}, /* 0xb5ac */
            {8'h00}, /* 0xb5ab */
            {8'h00}, /* 0xb5aa */
            {8'h00}, /* 0xb5a9 */
            {8'h00}, /* 0xb5a8 */
            {8'h00}, /* 0xb5a7 */
            {8'h00}, /* 0xb5a6 */
            {8'h00}, /* 0xb5a5 */
            {8'h00}, /* 0xb5a4 */
            {8'h00}, /* 0xb5a3 */
            {8'h00}, /* 0xb5a2 */
            {8'h00}, /* 0xb5a1 */
            {8'h00}, /* 0xb5a0 */
            {8'h00}, /* 0xb59f */
            {8'h00}, /* 0xb59e */
            {8'h00}, /* 0xb59d */
            {8'h00}, /* 0xb59c */
            {8'h00}, /* 0xb59b */
            {8'h00}, /* 0xb59a */
            {8'h00}, /* 0xb599 */
            {8'h00}, /* 0xb598 */
            {8'h00}, /* 0xb597 */
            {8'h00}, /* 0xb596 */
            {8'h00}, /* 0xb595 */
            {8'h00}, /* 0xb594 */
            {8'h00}, /* 0xb593 */
            {8'h00}, /* 0xb592 */
            {8'h00}, /* 0xb591 */
            {8'h00}, /* 0xb590 */
            {8'h00}, /* 0xb58f */
            {8'h00}, /* 0xb58e */
            {8'h00}, /* 0xb58d */
            {8'h00}, /* 0xb58c */
            {8'h00}, /* 0xb58b */
            {8'h00}, /* 0xb58a */
            {8'h00}, /* 0xb589 */
            {8'h00}, /* 0xb588 */
            {8'h00}, /* 0xb587 */
            {8'h00}, /* 0xb586 */
            {8'h00}, /* 0xb585 */
            {8'h00}, /* 0xb584 */
            {8'h00}, /* 0xb583 */
            {8'h00}, /* 0xb582 */
            {8'h00}, /* 0xb581 */
            {8'h00}, /* 0xb580 */
            {8'h00}, /* 0xb57f */
            {8'h00}, /* 0xb57e */
            {8'h00}, /* 0xb57d */
            {8'h00}, /* 0xb57c */
            {8'h00}, /* 0xb57b */
            {8'h00}, /* 0xb57a */
            {8'h00}, /* 0xb579 */
            {8'h00}, /* 0xb578 */
            {8'h00}, /* 0xb577 */
            {8'h00}, /* 0xb576 */
            {8'h00}, /* 0xb575 */
            {8'h00}, /* 0xb574 */
            {8'h00}, /* 0xb573 */
            {8'h00}, /* 0xb572 */
            {8'h00}, /* 0xb571 */
            {8'h00}, /* 0xb570 */
            {8'h00}, /* 0xb56f */
            {8'h00}, /* 0xb56e */
            {8'h00}, /* 0xb56d */
            {8'h00}, /* 0xb56c */
            {8'h00}, /* 0xb56b */
            {8'h00}, /* 0xb56a */
            {8'h00}, /* 0xb569 */
            {8'h00}, /* 0xb568 */
            {8'h00}, /* 0xb567 */
            {8'h00}, /* 0xb566 */
            {8'h00}, /* 0xb565 */
            {8'h00}, /* 0xb564 */
            {8'h00}, /* 0xb563 */
            {8'h00}, /* 0xb562 */
            {8'h00}, /* 0xb561 */
            {8'h00}, /* 0xb560 */
            {8'h00}, /* 0xb55f */
            {8'h00}, /* 0xb55e */
            {8'h00}, /* 0xb55d */
            {8'h00}, /* 0xb55c */
            {8'h00}, /* 0xb55b */
            {8'h00}, /* 0xb55a */
            {8'h00}, /* 0xb559 */
            {8'h00}, /* 0xb558 */
            {8'h00}, /* 0xb557 */
            {8'h00}, /* 0xb556 */
            {8'h00}, /* 0xb555 */
            {8'h00}, /* 0xb554 */
            {8'h00}, /* 0xb553 */
            {8'h00}, /* 0xb552 */
            {8'h00}, /* 0xb551 */
            {8'h00}, /* 0xb550 */
            {8'h00}, /* 0xb54f */
            {8'h00}, /* 0xb54e */
            {8'h00}, /* 0xb54d */
            {8'h00}, /* 0xb54c */
            {8'h00}, /* 0xb54b */
            {8'h00}, /* 0xb54a */
            {8'h00}, /* 0xb549 */
            {8'h00}, /* 0xb548 */
            {8'h00}, /* 0xb547 */
            {8'h00}, /* 0xb546 */
            {8'h00}, /* 0xb545 */
            {8'h00}, /* 0xb544 */
            {8'h00}, /* 0xb543 */
            {8'h00}, /* 0xb542 */
            {8'h00}, /* 0xb541 */
            {8'h00}, /* 0xb540 */
            {8'h00}, /* 0xb53f */
            {8'h00}, /* 0xb53e */
            {8'h00}, /* 0xb53d */
            {8'h00}, /* 0xb53c */
            {8'h00}, /* 0xb53b */
            {8'h00}, /* 0xb53a */
            {8'h00}, /* 0xb539 */
            {8'h00}, /* 0xb538 */
            {8'h00}, /* 0xb537 */
            {8'h00}, /* 0xb536 */
            {8'h00}, /* 0xb535 */
            {8'h00}, /* 0xb534 */
            {8'h00}, /* 0xb533 */
            {8'h00}, /* 0xb532 */
            {8'h00}, /* 0xb531 */
            {8'h00}, /* 0xb530 */
            {8'h00}, /* 0xb52f */
            {8'h00}, /* 0xb52e */
            {8'h00}, /* 0xb52d */
            {8'h00}, /* 0xb52c */
            {8'h00}, /* 0xb52b */
            {8'h00}, /* 0xb52a */
            {8'h00}, /* 0xb529 */
            {8'h00}, /* 0xb528 */
            {8'h00}, /* 0xb527 */
            {8'h00}, /* 0xb526 */
            {8'h00}, /* 0xb525 */
            {8'h00}, /* 0xb524 */
            {8'h00}, /* 0xb523 */
            {8'h00}, /* 0xb522 */
            {8'h00}, /* 0xb521 */
            {8'h00}, /* 0xb520 */
            {8'h00}, /* 0xb51f */
            {8'h00}, /* 0xb51e */
            {8'h00}, /* 0xb51d */
            {8'h00}, /* 0xb51c */
            {8'h00}, /* 0xb51b */
            {8'h00}, /* 0xb51a */
            {8'h00}, /* 0xb519 */
            {8'h00}, /* 0xb518 */
            {8'h00}, /* 0xb517 */
            {8'h00}, /* 0xb516 */
            {8'h00}, /* 0xb515 */
            {8'h00}, /* 0xb514 */
            {8'h00}, /* 0xb513 */
            {8'h00}, /* 0xb512 */
            {8'h00}, /* 0xb511 */
            {8'h00}, /* 0xb510 */
            {8'h00}, /* 0xb50f */
            {8'h00}, /* 0xb50e */
            {8'h00}, /* 0xb50d */
            {8'h00}, /* 0xb50c */
            {8'h00}, /* 0xb50b */
            {8'h00}, /* 0xb50a */
            {8'h00}, /* 0xb509 */
            {8'h00}, /* 0xb508 */
            {8'h00}, /* 0xb507 */
            {8'h00}, /* 0xb506 */
            {8'h00}, /* 0xb505 */
            {8'h00}, /* 0xb504 */
            {8'h00}, /* 0xb503 */
            {8'h00}, /* 0xb502 */
            {8'h00}, /* 0xb501 */
            {8'h00}, /* 0xb500 */
            {8'h00}, /* 0xb4ff */
            {8'h00}, /* 0xb4fe */
            {8'h00}, /* 0xb4fd */
            {8'h00}, /* 0xb4fc */
            {8'h00}, /* 0xb4fb */
            {8'h00}, /* 0xb4fa */
            {8'h00}, /* 0xb4f9 */
            {8'h00}, /* 0xb4f8 */
            {8'h00}, /* 0xb4f7 */
            {8'h00}, /* 0xb4f6 */
            {8'h00}, /* 0xb4f5 */
            {8'h00}, /* 0xb4f4 */
            {8'h00}, /* 0xb4f3 */
            {8'h00}, /* 0xb4f2 */
            {8'h00}, /* 0xb4f1 */
            {8'h00}, /* 0xb4f0 */
            {8'h00}, /* 0xb4ef */
            {8'h00}, /* 0xb4ee */
            {8'h00}, /* 0xb4ed */
            {8'h00}, /* 0xb4ec */
            {8'h00}, /* 0xb4eb */
            {8'h00}, /* 0xb4ea */
            {8'h00}, /* 0xb4e9 */
            {8'h00}, /* 0xb4e8 */
            {8'h00}, /* 0xb4e7 */
            {8'h00}, /* 0xb4e6 */
            {8'h00}, /* 0xb4e5 */
            {8'h00}, /* 0xb4e4 */
            {8'h00}, /* 0xb4e3 */
            {8'h00}, /* 0xb4e2 */
            {8'h00}, /* 0xb4e1 */
            {8'h00}, /* 0xb4e0 */
            {8'h00}, /* 0xb4df */
            {8'h00}, /* 0xb4de */
            {8'h00}, /* 0xb4dd */
            {8'h00}, /* 0xb4dc */
            {8'h00}, /* 0xb4db */
            {8'h00}, /* 0xb4da */
            {8'h00}, /* 0xb4d9 */
            {8'h00}, /* 0xb4d8 */
            {8'h00}, /* 0xb4d7 */
            {8'h00}, /* 0xb4d6 */
            {8'h00}, /* 0xb4d5 */
            {8'h00}, /* 0xb4d4 */
            {8'h00}, /* 0xb4d3 */
            {8'h00}, /* 0xb4d2 */
            {8'h00}, /* 0xb4d1 */
            {8'h00}, /* 0xb4d0 */
            {8'h00}, /* 0xb4cf */
            {8'h00}, /* 0xb4ce */
            {8'h00}, /* 0xb4cd */
            {8'h00}, /* 0xb4cc */
            {8'h00}, /* 0xb4cb */
            {8'h00}, /* 0xb4ca */
            {8'h00}, /* 0xb4c9 */
            {8'h00}, /* 0xb4c8 */
            {8'h00}, /* 0xb4c7 */
            {8'h00}, /* 0xb4c6 */
            {8'h00}, /* 0xb4c5 */
            {8'h00}, /* 0xb4c4 */
            {8'h00}, /* 0xb4c3 */
            {8'h00}, /* 0xb4c2 */
            {8'h00}, /* 0xb4c1 */
            {8'h00}, /* 0xb4c0 */
            {8'h00}, /* 0xb4bf */
            {8'h00}, /* 0xb4be */
            {8'h00}, /* 0xb4bd */
            {8'h00}, /* 0xb4bc */
            {8'h00}, /* 0xb4bb */
            {8'h00}, /* 0xb4ba */
            {8'h00}, /* 0xb4b9 */
            {8'h00}, /* 0xb4b8 */
            {8'h00}, /* 0xb4b7 */
            {8'h00}, /* 0xb4b6 */
            {8'h00}, /* 0xb4b5 */
            {8'h00}, /* 0xb4b4 */
            {8'h00}, /* 0xb4b3 */
            {8'h00}, /* 0xb4b2 */
            {8'h00}, /* 0xb4b1 */
            {8'h00}, /* 0xb4b0 */
            {8'h00}, /* 0xb4af */
            {8'h00}, /* 0xb4ae */
            {8'h00}, /* 0xb4ad */
            {8'h00}, /* 0xb4ac */
            {8'h00}, /* 0xb4ab */
            {8'h00}, /* 0xb4aa */
            {8'h00}, /* 0xb4a9 */
            {8'h00}, /* 0xb4a8 */
            {8'h00}, /* 0xb4a7 */
            {8'h00}, /* 0xb4a6 */
            {8'h00}, /* 0xb4a5 */
            {8'h00}, /* 0xb4a4 */
            {8'h00}, /* 0xb4a3 */
            {8'h00}, /* 0xb4a2 */
            {8'h00}, /* 0xb4a1 */
            {8'h00}, /* 0xb4a0 */
            {8'h00}, /* 0xb49f */
            {8'h00}, /* 0xb49e */
            {8'h00}, /* 0xb49d */
            {8'h00}, /* 0xb49c */
            {8'h00}, /* 0xb49b */
            {8'h00}, /* 0xb49a */
            {8'h00}, /* 0xb499 */
            {8'h00}, /* 0xb498 */
            {8'h00}, /* 0xb497 */
            {8'h00}, /* 0xb496 */
            {8'h00}, /* 0xb495 */
            {8'h00}, /* 0xb494 */
            {8'h00}, /* 0xb493 */
            {8'h00}, /* 0xb492 */
            {8'h00}, /* 0xb491 */
            {8'h00}, /* 0xb490 */
            {8'h00}, /* 0xb48f */
            {8'h00}, /* 0xb48e */
            {8'h00}, /* 0xb48d */
            {8'h00}, /* 0xb48c */
            {8'h00}, /* 0xb48b */
            {8'h00}, /* 0xb48a */
            {8'h00}, /* 0xb489 */
            {8'h00}, /* 0xb488 */
            {8'h00}, /* 0xb487 */
            {8'h00}, /* 0xb486 */
            {8'h00}, /* 0xb485 */
            {8'h00}, /* 0xb484 */
            {8'h00}, /* 0xb483 */
            {8'h00}, /* 0xb482 */
            {8'h00}, /* 0xb481 */
            {8'h00}, /* 0xb480 */
            {8'h00}, /* 0xb47f */
            {8'h00}, /* 0xb47e */
            {8'h00}, /* 0xb47d */
            {8'h00}, /* 0xb47c */
            {8'h00}, /* 0xb47b */
            {8'h00}, /* 0xb47a */
            {8'h00}, /* 0xb479 */
            {8'h00}, /* 0xb478 */
            {8'h00}, /* 0xb477 */
            {8'h00}, /* 0xb476 */
            {8'h00}, /* 0xb475 */
            {8'h00}, /* 0xb474 */
            {8'h00}, /* 0xb473 */
            {8'h00}, /* 0xb472 */
            {8'h00}, /* 0xb471 */
            {8'h00}, /* 0xb470 */
            {8'h00}, /* 0xb46f */
            {8'h00}, /* 0xb46e */
            {8'h00}, /* 0xb46d */
            {8'h00}, /* 0xb46c */
            {8'h00}, /* 0xb46b */
            {8'h00}, /* 0xb46a */
            {8'h00}, /* 0xb469 */
            {8'h00}, /* 0xb468 */
            {8'h00}, /* 0xb467 */
            {8'h00}, /* 0xb466 */
            {8'h00}, /* 0xb465 */
            {8'h00}, /* 0xb464 */
            {8'h00}, /* 0xb463 */
            {8'h00}, /* 0xb462 */
            {8'h00}, /* 0xb461 */
            {8'h00}, /* 0xb460 */
            {8'h00}, /* 0xb45f */
            {8'h00}, /* 0xb45e */
            {8'h00}, /* 0xb45d */
            {8'h00}, /* 0xb45c */
            {8'h00}, /* 0xb45b */
            {8'h00}, /* 0xb45a */
            {8'h00}, /* 0xb459 */
            {8'h00}, /* 0xb458 */
            {8'h00}, /* 0xb457 */
            {8'h00}, /* 0xb456 */
            {8'h00}, /* 0xb455 */
            {8'h00}, /* 0xb454 */
            {8'h00}, /* 0xb453 */
            {8'h00}, /* 0xb452 */
            {8'h00}, /* 0xb451 */
            {8'h00}, /* 0xb450 */
            {8'h00}, /* 0xb44f */
            {8'h00}, /* 0xb44e */
            {8'h00}, /* 0xb44d */
            {8'h00}, /* 0xb44c */
            {8'h00}, /* 0xb44b */
            {8'h00}, /* 0xb44a */
            {8'h00}, /* 0xb449 */
            {8'h00}, /* 0xb448 */
            {8'h00}, /* 0xb447 */
            {8'h00}, /* 0xb446 */
            {8'h00}, /* 0xb445 */
            {8'h00}, /* 0xb444 */
            {8'h00}, /* 0xb443 */
            {8'h00}, /* 0xb442 */
            {8'h00}, /* 0xb441 */
            {8'h00}, /* 0xb440 */
            {8'h00}, /* 0xb43f */
            {8'h00}, /* 0xb43e */
            {8'h00}, /* 0xb43d */
            {8'h00}, /* 0xb43c */
            {8'h00}, /* 0xb43b */
            {8'h00}, /* 0xb43a */
            {8'h00}, /* 0xb439 */
            {8'h00}, /* 0xb438 */
            {8'h00}, /* 0xb437 */
            {8'h00}, /* 0xb436 */
            {8'h00}, /* 0xb435 */
            {8'h00}, /* 0xb434 */
            {8'h00}, /* 0xb433 */
            {8'h00}, /* 0xb432 */
            {8'h00}, /* 0xb431 */
            {8'h00}, /* 0xb430 */
            {8'h00}, /* 0xb42f */
            {8'h00}, /* 0xb42e */
            {8'h00}, /* 0xb42d */
            {8'h00}, /* 0xb42c */
            {8'h00}, /* 0xb42b */
            {8'h00}, /* 0xb42a */
            {8'h00}, /* 0xb429 */
            {8'h00}, /* 0xb428 */
            {8'h00}, /* 0xb427 */
            {8'h00}, /* 0xb426 */
            {8'h00}, /* 0xb425 */
            {8'h00}, /* 0xb424 */
            {8'h00}, /* 0xb423 */
            {8'h00}, /* 0xb422 */
            {8'h00}, /* 0xb421 */
            {8'h00}, /* 0xb420 */
            {8'h00}, /* 0xb41f */
            {8'h00}, /* 0xb41e */
            {8'h00}, /* 0xb41d */
            {8'h00}, /* 0xb41c */
            {8'h00}, /* 0xb41b */
            {8'h00}, /* 0xb41a */
            {8'h00}, /* 0xb419 */
            {8'h00}, /* 0xb418 */
            {8'h00}, /* 0xb417 */
            {8'h00}, /* 0xb416 */
            {8'h00}, /* 0xb415 */
            {8'h00}, /* 0xb414 */
            {8'h00}, /* 0xb413 */
            {8'h00}, /* 0xb412 */
            {8'h00}, /* 0xb411 */
            {8'h00}, /* 0xb410 */
            {8'h00}, /* 0xb40f */
            {8'h00}, /* 0xb40e */
            {8'h00}, /* 0xb40d */
            {8'h00}, /* 0xb40c */
            {8'h00}, /* 0xb40b */
            {8'h00}, /* 0xb40a */
            {8'h00}, /* 0xb409 */
            {8'h00}, /* 0xb408 */
            {8'h00}, /* 0xb407 */
            {8'h00}, /* 0xb406 */
            {8'h00}, /* 0xb405 */
            {8'h00}, /* 0xb404 */
            {8'h00}, /* 0xb403 */
            {8'h00}, /* 0xb402 */
            {8'h00}, /* 0xb401 */
            {8'h00}, /* 0xb400 */
            {8'h00}, /* 0xb3ff */
            {8'h00}, /* 0xb3fe */
            {8'h00}, /* 0xb3fd */
            {8'h00}, /* 0xb3fc */
            {8'h00}, /* 0xb3fb */
            {8'h00}, /* 0xb3fa */
            {8'h00}, /* 0xb3f9 */
            {8'h00}, /* 0xb3f8 */
            {8'h00}, /* 0xb3f7 */
            {8'h00}, /* 0xb3f6 */
            {8'h00}, /* 0xb3f5 */
            {8'h00}, /* 0xb3f4 */
            {8'h00}, /* 0xb3f3 */
            {8'h00}, /* 0xb3f2 */
            {8'h00}, /* 0xb3f1 */
            {8'h00}, /* 0xb3f0 */
            {8'h00}, /* 0xb3ef */
            {8'h00}, /* 0xb3ee */
            {8'h00}, /* 0xb3ed */
            {8'h00}, /* 0xb3ec */
            {8'h00}, /* 0xb3eb */
            {8'h00}, /* 0xb3ea */
            {8'h00}, /* 0xb3e9 */
            {8'h00}, /* 0xb3e8 */
            {8'h00}, /* 0xb3e7 */
            {8'h00}, /* 0xb3e6 */
            {8'h00}, /* 0xb3e5 */
            {8'h00}, /* 0xb3e4 */
            {8'h00}, /* 0xb3e3 */
            {8'h00}, /* 0xb3e2 */
            {8'h00}, /* 0xb3e1 */
            {8'h00}, /* 0xb3e0 */
            {8'h00}, /* 0xb3df */
            {8'h00}, /* 0xb3de */
            {8'h00}, /* 0xb3dd */
            {8'h00}, /* 0xb3dc */
            {8'h00}, /* 0xb3db */
            {8'h00}, /* 0xb3da */
            {8'h00}, /* 0xb3d9 */
            {8'h00}, /* 0xb3d8 */
            {8'h00}, /* 0xb3d7 */
            {8'h00}, /* 0xb3d6 */
            {8'h00}, /* 0xb3d5 */
            {8'h00}, /* 0xb3d4 */
            {8'h00}, /* 0xb3d3 */
            {8'h00}, /* 0xb3d2 */
            {8'h00}, /* 0xb3d1 */
            {8'h00}, /* 0xb3d0 */
            {8'h00}, /* 0xb3cf */
            {8'h00}, /* 0xb3ce */
            {8'h00}, /* 0xb3cd */
            {8'h00}, /* 0xb3cc */
            {8'h00}, /* 0xb3cb */
            {8'h00}, /* 0xb3ca */
            {8'h00}, /* 0xb3c9 */
            {8'h00}, /* 0xb3c8 */
            {8'h00}, /* 0xb3c7 */
            {8'h00}, /* 0xb3c6 */
            {8'h00}, /* 0xb3c5 */
            {8'h00}, /* 0xb3c4 */
            {8'h00}, /* 0xb3c3 */
            {8'h00}, /* 0xb3c2 */
            {8'h00}, /* 0xb3c1 */
            {8'h00}, /* 0xb3c0 */
            {8'h00}, /* 0xb3bf */
            {8'h00}, /* 0xb3be */
            {8'h00}, /* 0xb3bd */
            {8'h00}, /* 0xb3bc */
            {8'h00}, /* 0xb3bb */
            {8'h00}, /* 0xb3ba */
            {8'h00}, /* 0xb3b9 */
            {8'h00}, /* 0xb3b8 */
            {8'h00}, /* 0xb3b7 */
            {8'h00}, /* 0xb3b6 */
            {8'h00}, /* 0xb3b5 */
            {8'h00}, /* 0xb3b4 */
            {8'h00}, /* 0xb3b3 */
            {8'h00}, /* 0xb3b2 */
            {8'h00}, /* 0xb3b1 */
            {8'h00}, /* 0xb3b0 */
            {8'h00}, /* 0xb3af */
            {8'h00}, /* 0xb3ae */
            {8'h00}, /* 0xb3ad */
            {8'h00}, /* 0xb3ac */
            {8'h00}, /* 0xb3ab */
            {8'h00}, /* 0xb3aa */
            {8'h00}, /* 0xb3a9 */
            {8'h00}, /* 0xb3a8 */
            {8'h00}, /* 0xb3a7 */
            {8'h00}, /* 0xb3a6 */
            {8'h00}, /* 0xb3a5 */
            {8'h00}, /* 0xb3a4 */
            {8'h00}, /* 0xb3a3 */
            {8'h00}, /* 0xb3a2 */
            {8'h00}, /* 0xb3a1 */
            {8'h00}, /* 0xb3a0 */
            {8'h00}, /* 0xb39f */
            {8'h00}, /* 0xb39e */
            {8'h00}, /* 0xb39d */
            {8'h00}, /* 0xb39c */
            {8'h00}, /* 0xb39b */
            {8'h00}, /* 0xb39a */
            {8'h00}, /* 0xb399 */
            {8'h00}, /* 0xb398 */
            {8'h00}, /* 0xb397 */
            {8'h00}, /* 0xb396 */
            {8'h00}, /* 0xb395 */
            {8'h00}, /* 0xb394 */
            {8'h00}, /* 0xb393 */
            {8'h00}, /* 0xb392 */
            {8'h00}, /* 0xb391 */
            {8'h00}, /* 0xb390 */
            {8'h00}, /* 0xb38f */
            {8'h00}, /* 0xb38e */
            {8'h00}, /* 0xb38d */
            {8'h00}, /* 0xb38c */
            {8'h00}, /* 0xb38b */
            {8'h00}, /* 0xb38a */
            {8'h00}, /* 0xb389 */
            {8'h00}, /* 0xb388 */
            {8'h00}, /* 0xb387 */
            {8'h00}, /* 0xb386 */
            {8'h00}, /* 0xb385 */
            {8'h00}, /* 0xb384 */
            {8'h00}, /* 0xb383 */
            {8'h00}, /* 0xb382 */
            {8'h00}, /* 0xb381 */
            {8'h00}, /* 0xb380 */
            {8'h00}, /* 0xb37f */
            {8'h00}, /* 0xb37e */
            {8'h00}, /* 0xb37d */
            {8'h00}, /* 0xb37c */
            {8'h00}, /* 0xb37b */
            {8'h00}, /* 0xb37a */
            {8'h00}, /* 0xb379 */
            {8'h00}, /* 0xb378 */
            {8'h00}, /* 0xb377 */
            {8'h00}, /* 0xb376 */
            {8'h00}, /* 0xb375 */
            {8'h00}, /* 0xb374 */
            {8'h00}, /* 0xb373 */
            {8'h00}, /* 0xb372 */
            {8'h00}, /* 0xb371 */
            {8'h00}, /* 0xb370 */
            {8'h00}, /* 0xb36f */
            {8'h00}, /* 0xb36e */
            {8'h00}, /* 0xb36d */
            {8'h00}, /* 0xb36c */
            {8'h00}, /* 0xb36b */
            {8'h00}, /* 0xb36a */
            {8'h00}, /* 0xb369 */
            {8'h00}, /* 0xb368 */
            {8'h00}, /* 0xb367 */
            {8'h00}, /* 0xb366 */
            {8'h00}, /* 0xb365 */
            {8'h00}, /* 0xb364 */
            {8'h00}, /* 0xb363 */
            {8'h00}, /* 0xb362 */
            {8'h00}, /* 0xb361 */
            {8'h00}, /* 0xb360 */
            {8'h00}, /* 0xb35f */
            {8'h00}, /* 0xb35e */
            {8'h00}, /* 0xb35d */
            {8'h00}, /* 0xb35c */
            {8'h00}, /* 0xb35b */
            {8'h00}, /* 0xb35a */
            {8'h00}, /* 0xb359 */
            {8'h00}, /* 0xb358 */
            {8'h00}, /* 0xb357 */
            {8'h00}, /* 0xb356 */
            {8'h00}, /* 0xb355 */
            {8'h00}, /* 0xb354 */
            {8'h00}, /* 0xb353 */
            {8'h00}, /* 0xb352 */
            {8'h00}, /* 0xb351 */
            {8'h00}, /* 0xb350 */
            {8'h00}, /* 0xb34f */
            {8'h00}, /* 0xb34e */
            {8'h00}, /* 0xb34d */
            {8'h00}, /* 0xb34c */
            {8'h00}, /* 0xb34b */
            {8'h00}, /* 0xb34a */
            {8'h00}, /* 0xb349 */
            {8'h00}, /* 0xb348 */
            {8'h00}, /* 0xb347 */
            {8'h00}, /* 0xb346 */
            {8'h00}, /* 0xb345 */
            {8'h00}, /* 0xb344 */
            {8'h00}, /* 0xb343 */
            {8'h00}, /* 0xb342 */
            {8'h00}, /* 0xb341 */
            {8'h00}, /* 0xb340 */
            {8'h00}, /* 0xb33f */
            {8'h00}, /* 0xb33e */
            {8'h00}, /* 0xb33d */
            {8'h00}, /* 0xb33c */
            {8'h00}, /* 0xb33b */
            {8'h00}, /* 0xb33a */
            {8'h00}, /* 0xb339 */
            {8'h00}, /* 0xb338 */
            {8'h00}, /* 0xb337 */
            {8'h00}, /* 0xb336 */
            {8'h00}, /* 0xb335 */
            {8'h00}, /* 0xb334 */
            {8'h00}, /* 0xb333 */
            {8'h00}, /* 0xb332 */
            {8'h00}, /* 0xb331 */
            {8'h00}, /* 0xb330 */
            {8'h00}, /* 0xb32f */
            {8'h00}, /* 0xb32e */
            {8'h00}, /* 0xb32d */
            {8'h00}, /* 0xb32c */
            {8'h00}, /* 0xb32b */
            {8'h00}, /* 0xb32a */
            {8'h00}, /* 0xb329 */
            {8'h00}, /* 0xb328 */
            {8'h00}, /* 0xb327 */
            {8'h00}, /* 0xb326 */
            {8'h00}, /* 0xb325 */
            {8'h00}, /* 0xb324 */
            {8'h00}, /* 0xb323 */
            {8'h00}, /* 0xb322 */
            {8'h00}, /* 0xb321 */
            {8'h00}, /* 0xb320 */
            {8'h00}, /* 0xb31f */
            {8'h00}, /* 0xb31e */
            {8'h00}, /* 0xb31d */
            {8'h00}, /* 0xb31c */
            {8'h00}, /* 0xb31b */
            {8'h00}, /* 0xb31a */
            {8'h00}, /* 0xb319 */
            {8'h00}, /* 0xb318 */
            {8'h00}, /* 0xb317 */
            {8'h00}, /* 0xb316 */
            {8'h00}, /* 0xb315 */
            {8'h00}, /* 0xb314 */
            {8'h00}, /* 0xb313 */
            {8'h00}, /* 0xb312 */
            {8'h00}, /* 0xb311 */
            {8'h00}, /* 0xb310 */
            {8'h00}, /* 0xb30f */
            {8'h00}, /* 0xb30e */
            {8'h00}, /* 0xb30d */
            {8'h00}, /* 0xb30c */
            {8'h00}, /* 0xb30b */
            {8'h00}, /* 0xb30a */
            {8'h00}, /* 0xb309 */
            {8'h00}, /* 0xb308 */
            {8'h00}, /* 0xb307 */
            {8'h00}, /* 0xb306 */
            {8'h00}, /* 0xb305 */
            {8'h00}, /* 0xb304 */
            {8'h00}, /* 0xb303 */
            {8'h00}, /* 0xb302 */
            {8'h00}, /* 0xb301 */
            {8'h00}, /* 0xb300 */
            {8'h00}, /* 0xb2ff */
            {8'h00}, /* 0xb2fe */
            {8'h00}, /* 0xb2fd */
            {8'h00}, /* 0xb2fc */
            {8'h00}, /* 0xb2fb */
            {8'h00}, /* 0xb2fa */
            {8'h00}, /* 0xb2f9 */
            {8'h00}, /* 0xb2f8 */
            {8'h00}, /* 0xb2f7 */
            {8'h00}, /* 0xb2f6 */
            {8'h00}, /* 0xb2f5 */
            {8'h00}, /* 0xb2f4 */
            {8'h00}, /* 0xb2f3 */
            {8'h00}, /* 0xb2f2 */
            {8'h00}, /* 0xb2f1 */
            {8'h00}, /* 0xb2f0 */
            {8'h00}, /* 0xb2ef */
            {8'h00}, /* 0xb2ee */
            {8'h00}, /* 0xb2ed */
            {8'h00}, /* 0xb2ec */
            {8'h00}, /* 0xb2eb */
            {8'h00}, /* 0xb2ea */
            {8'h00}, /* 0xb2e9 */
            {8'h00}, /* 0xb2e8 */
            {8'h00}, /* 0xb2e7 */
            {8'h00}, /* 0xb2e6 */
            {8'h00}, /* 0xb2e5 */
            {8'h00}, /* 0xb2e4 */
            {8'h00}, /* 0xb2e3 */
            {8'h00}, /* 0xb2e2 */
            {8'h00}, /* 0xb2e1 */
            {8'h00}, /* 0xb2e0 */
            {8'h00}, /* 0xb2df */
            {8'h00}, /* 0xb2de */
            {8'h00}, /* 0xb2dd */
            {8'h00}, /* 0xb2dc */
            {8'h00}, /* 0xb2db */
            {8'h00}, /* 0xb2da */
            {8'h00}, /* 0xb2d9 */
            {8'h00}, /* 0xb2d8 */
            {8'h00}, /* 0xb2d7 */
            {8'h00}, /* 0xb2d6 */
            {8'h00}, /* 0xb2d5 */
            {8'h00}, /* 0xb2d4 */
            {8'h00}, /* 0xb2d3 */
            {8'h00}, /* 0xb2d2 */
            {8'h00}, /* 0xb2d1 */
            {8'h00}, /* 0xb2d0 */
            {8'h00}, /* 0xb2cf */
            {8'h00}, /* 0xb2ce */
            {8'h00}, /* 0xb2cd */
            {8'h00}, /* 0xb2cc */
            {8'h00}, /* 0xb2cb */
            {8'h00}, /* 0xb2ca */
            {8'h00}, /* 0xb2c9 */
            {8'h00}, /* 0xb2c8 */
            {8'h00}, /* 0xb2c7 */
            {8'h00}, /* 0xb2c6 */
            {8'h00}, /* 0xb2c5 */
            {8'h00}, /* 0xb2c4 */
            {8'h00}, /* 0xb2c3 */
            {8'h00}, /* 0xb2c2 */
            {8'h00}, /* 0xb2c1 */
            {8'h00}, /* 0xb2c0 */
            {8'h00}, /* 0xb2bf */
            {8'h00}, /* 0xb2be */
            {8'h00}, /* 0xb2bd */
            {8'h00}, /* 0xb2bc */
            {8'h00}, /* 0xb2bb */
            {8'h00}, /* 0xb2ba */
            {8'h00}, /* 0xb2b9 */
            {8'h00}, /* 0xb2b8 */
            {8'h00}, /* 0xb2b7 */
            {8'h00}, /* 0xb2b6 */
            {8'h00}, /* 0xb2b5 */
            {8'h00}, /* 0xb2b4 */
            {8'h00}, /* 0xb2b3 */
            {8'h00}, /* 0xb2b2 */
            {8'h00}, /* 0xb2b1 */
            {8'h00}, /* 0xb2b0 */
            {8'h00}, /* 0xb2af */
            {8'h00}, /* 0xb2ae */
            {8'h00}, /* 0xb2ad */
            {8'h00}, /* 0xb2ac */
            {8'h00}, /* 0xb2ab */
            {8'h00}, /* 0xb2aa */
            {8'h00}, /* 0xb2a9 */
            {8'h00}, /* 0xb2a8 */
            {8'h00}, /* 0xb2a7 */
            {8'h00}, /* 0xb2a6 */
            {8'h00}, /* 0xb2a5 */
            {8'h00}, /* 0xb2a4 */
            {8'h00}, /* 0xb2a3 */
            {8'h00}, /* 0xb2a2 */
            {8'h00}, /* 0xb2a1 */
            {8'h00}, /* 0xb2a0 */
            {8'h00}, /* 0xb29f */
            {8'h00}, /* 0xb29e */
            {8'h00}, /* 0xb29d */
            {8'h00}, /* 0xb29c */
            {8'h00}, /* 0xb29b */
            {8'h00}, /* 0xb29a */
            {8'h00}, /* 0xb299 */
            {8'h00}, /* 0xb298 */
            {8'h00}, /* 0xb297 */
            {8'h00}, /* 0xb296 */
            {8'h00}, /* 0xb295 */
            {8'h00}, /* 0xb294 */
            {8'h00}, /* 0xb293 */
            {8'h00}, /* 0xb292 */
            {8'h00}, /* 0xb291 */
            {8'h00}, /* 0xb290 */
            {8'h00}, /* 0xb28f */
            {8'h00}, /* 0xb28e */
            {8'h00}, /* 0xb28d */
            {8'h00}, /* 0xb28c */
            {8'h00}, /* 0xb28b */
            {8'h00}, /* 0xb28a */
            {8'h00}, /* 0xb289 */
            {8'h00}, /* 0xb288 */
            {8'h00}, /* 0xb287 */
            {8'h00}, /* 0xb286 */
            {8'h00}, /* 0xb285 */
            {8'h00}, /* 0xb284 */
            {8'h00}, /* 0xb283 */
            {8'h00}, /* 0xb282 */
            {8'h00}, /* 0xb281 */
            {8'h00}, /* 0xb280 */
            {8'h00}, /* 0xb27f */
            {8'h00}, /* 0xb27e */
            {8'h00}, /* 0xb27d */
            {8'h00}, /* 0xb27c */
            {8'h00}, /* 0xb27b */
            {8'h00}, /* 0xb27a */
            {8'h00}, /* 0xb279 */
            {8'h00}, /* 0xb278 */
            {8'h00}, /* 0xb277 */
            {8'h00}, /* 0xb276 */
            {8'h00}, /* 0xb275 */
            {8'h00}, /* 0xb274 */
            {8'h00}, /* 0xb273 */
            {8'h00}, /* 0xb272 */
            {8'h00}, /* 0xb271 */
            {8'h00}, /* 0xb270 */
            {8'h00}, /* 0xb26f */
            {8'h00}, /* 0xb26e */
            {8'h00}, /* 0xb26d */
            {8'h00}, /* 0xb26c */
            {8'h00}, /* 0xb26b */
            {8'h00}, /* 0xb26a */
            {8'h00}, /* 0xb269 */
            {8'h00}, /* 0xb268 */
            {8'h00}, /* 0xb267 */
            {8'h00}, /* 0xb266 */
            {8'h00}, /* 0xb265 */
            {8'h00}, /* 0xb264 */
            {8'h00}, /* 0xb263 */
            {8'h00}, /* 0xb262 */
            {8'h00}, /* 0xb261 */
            {8'h00}, /* 0xb260 */
            {8'h00}, /* 0xb25f */
            {8'h00}, /* 0xb25e */
            {8'h00}, /* 0xb25d */
            {8'h00}, /* 0xb25c */
            {8'h00}, /* 0xb25b */
            {8'h00}, /* 0xb25a */
            {8'h00}, /* 0xb259 */
            {8'h00}, /* 0xb258 */
            {8'h00}, /* 0xb257 */
            {8'h00}, /* 0xb256 */
            {8'h00}, /* 0xb255 */
            {8'h00}, /* 0xb254 */
            {8'h00}, /* 0xb253 */
            {8'h00}, /* 0xb252 */
            {8'h00}, /* 0xb251 */
            {8'h00}, /* 0xb250 */
            {8'h00}, /* 0xb24f */
            {8'h00}, /* 0xb24e */
            {8'h00}, /* 0xb24d */
            {8'h00}, /* 0xb24c */
            {8'h00}, /* 0xb24b */
            {8'h00}, /* 0xb24a */
            {8'h00}, /* 0xb249 */
            {8'h00}, /* 0xb248 */
            {8'h00}, /* 0xb247 */
            {8'h00}, /* 0xb246 */
            {8'h00}, /* 0xb245 */
            {8'h00}, /* 0xb244 */
            {8'h00}, /* 0xb243 */
            {8'h00}, /* 0xb242 */
            {8'h00}, /* 0xb241 */
            {8'h00}, /* 0xb240 */
            {8'h00}, /* 0xb23f */
            {8'h00}, /* 0xb23e */
            {8'h00}, /* 0xb23d */
            {8'h00}, /* 0xb23c */
            {8'h00}, /* 0xb23b */
            {8'h00}, /* 0xb23a */
            {8'h00}, /* 0xb239 */
            {8'h00}, /* 0xb238 */
            {8'h00}, /* 0xb237 */
            {8'h00}, /* 0xb236 */
            {8'h00}, /* 0xb235 */
            {8'h00}, /* 0xb234 */
            {8'h00}, /* 0xb233 */
            {8'h00}, /* 0xb232 */
            {8'h00}, /* 0xb231 */
            {8'h00}, /* 0xb230 */
            {8'h00}, /* 0xb22f */
            {8'h00}, /* 0xb22e */
            {8'h00}, /* 0xb22d */
            {8'h00}, /* 0xb22c */
            {8'h00}, /* 0xb22b */
            {8'h00}, /* 0xb22a */
            {8'h00}, /* 0xb229 */
            {8'h00}, /* 0xb228 */
            {8'h00}, /* 0xb227 */
            {8'h00}, /* 0xb226 */
            {8'h00}, /* 0xb225 */
            {8'h00}, /* 0xb224 */
            {8'h00}, /* 0xb223 */
            {8'h00}, /* 0xb222 */
            {8'h00}, /* 0xb221 */
            {8'h00}, /* 0xb220 */
            {8'h00}, /* 0xb21f */
            {8'h00}, /* 0xb21e */
            {8'h00}, /* 0xb21d */
            {8'h00}, /* 0xb21c */
            {8'h00}, /* 0xb21b */
            {8'h00}, /* 0xb21a */
            {8'h00}, /* 0xb219 */
            {8'h00}, /* 0xb218 */
            {8'h00}, /* 0xb217 */
            {8'h00}, /* 0xb216 */
            {8'h00}, /* 0xb215 */
            {8'h00}, /* 0xb214 */
            {8'h00}, /* 0xb213 */
            {8'h00}, /* 0xb212 */
            {8'h00}, /* 0xb211 */
            {8'h00}, /* 0xb210 */
            {8'h00}, /* 0xb20f */
            {8'h00}, /* 0xb20e */
            {8'h00}, /* 0xb20d */
            {8'h00}, /* 0xb20c */
            {8'h00}, /* 0xb20b */
            {8'h00}, /* 0xb20a */
            {8'h00}, /* 0xb209 */
            {8'h00}, /* 0xb208 */
            {8'h00}, /* 0xb207 */
            {8'h00}, /* 0xb206 */
            {8'h00}, /* 0xb205 */
            {8'h00}, /* 0xb204 */
            {8'h00}, /* 0xb203 */
            {8'h00}, /* 0xb202 */
            {8'h00}, /* 0xb201 */
            {8'h00}, /* 0xb200 */
            {8'h00}, /* 0xb1ff */
            {8'h00}, /* 0xb1fe */
            {8'h00}, /* 0xb1fd */
            {8'h00}, /* 0xb1fc */
            {8'h00}, /* 0xb1fb */
            {8'h00}, /* 0xb1fa */
            {8'h00}, /* 0xb1f9 */
            {8'h00}, /* 0xb1f8 */
            {8'h00}, /* 0xb1f7 */
            {8'h00}, /* 0xb1f6 */
            {8'h00}, /* 0xb1f5 */
            {8'h00}, /* 0xb1f4 */
            {8'h00}, /* 0xb1f3 */
            {8'h00}, /* 0xb1f2 */
            {8'h00}, /* 0xb1f1 */
            {8'h00}, /* 0xb1f0 */
            {8'h00}, /* 0xb1ef */
            {8'h00}, /* 0xb1ee */
            {8'h00}, /* 0xb1ed */
            {8'h00}, /* 0xb1ec */
            {8'h00}, /* 0xb1eb */
            {8'h00}, /* 0xb1ea */
            {8'h00}, /* 0xb1e9 */
            {8'h00}, /* 0xb1e8 */
            {8'h00}, /* 0xb1e7 */
            {8'h00}, /* 0xb1e6 */
            {8'h00}, /* 0xb1e5 */
            {8'h00}, /* 0xb1e4 */
            {8'h00}, /* 0xb1e3 */
            {8'h00}, /* 0xb1e2 */
            {8'h00}, /* 0xb1e1 */
            {8'h00}, /* 0xb1e0 */
            {8'h00}, /* 0xb1df */
            {8'h00}, /* 0xb1de */
            {8'h00}, /* 0xb1dd */
            {8'h00}, /* 0xb1dc */
            {8'h00}, /* 0xb1db */
            {8'h00}, /* 0xb1da */
            {8'h00}, /* 0xb1d9 */
            {8'h00}, /* 0xb1d8 */
            {8'h00}, /* 0xb1d7 */
            {8'h00}, /* 0xb1d6 */
            {8'h00}, /* 0xb1d5 */
            {8'h00}, /* 0xb1d4 */
            {8'h00}, /* 0xb1d3 */
            {8'h00}, /* 0xb1d2 */
            {8'h00}, /* 0xb1d1 */
            {8'h00}, /* 0xb1d0 */
            {8'h00}, /* 0xb1cf */
            {8'h00}, /* 0xb1ce */
            {8'h00}, /* 0xb1cd */
            {8'h00}, /* 0xb1cc */
            {8'h00}, /* 0xb1cb */
            {8'h00}, /* 0xb1ca */
            {8'h00}, /* 0xb1c9 */
            {8'h00}, /* 0xb1c8 */
            {8'h00}, /* 0xb1c7 */
            {8'h00}, /* 0xb1c6 */
            {8'h00}, /* 0xb1c5 */
            {8'h00}, /* 0xb1c4 */
            {8'h00}, /* 0xb1c3 */
            {8'h00}, /* 0xb1c2 */
            {8'h00}, /* 0xb1c1 */
            {8'h00}, /* 0xb1c0 */
            {8'h00}, /* 0xb1bf */
            {8'h00}, /* 0xb1be */
            {8'h00}, /* 0xb1bd */
            {8'h00}, /* 0xb1bc */
            {8'h00}, /* 0xb1bb */
            {8'h00}, /* 0xb1ba */
            {8'h00}, /* 0xb1b9 */
            {8'h00}, /* 0xb1b8 */
            {8'h00}, /* 0xb1b7 */
            {8'h00}, /* 0xb1b6 */
            {8'h00}, /* 0xb1b5 */
            {8'h00}, /* 0xb1b4 */
            {8'h00}, /* 0xb1b3 */
            {8'h00}, /* 0xb1b2 */
            {8'h00}, /* 0xb1b1 */
            {8'h00}, /* 0xb1b0 */
            {8'h00}, /* 0xb1af */
            {8'h00}, /* 0xb1ae */
            {8'h00}, /* 0xb1ad */
            {8'h00}, /* 0xb1ac */
            {8'h00}, /* 0xb1ab */
            {8'h00}, /* 0xb1aa */
            {8'h00}, /* 0xb1a9 */
            {8'h00}, /* 0xb1a8 */
            {8'h00}, /* 0xb1a7 */
            {8'h00}, /* 0xb1a6 */
            {8'h00}, /* 0xb1a5 */
            {8'h00}, /* 0xb1a4 */
            {8'h00}, /* 0xb1a3 */
            {8'h00}, /* 0xb1a2 */
            {8'h00}, /* 0xb1a1 */
            {8'h00}, /* 0xb1a0 */
            {8'h00}, /* 0xb19f */
            {8'h00}, /* 0xb19e */
            {8'h00}, /* 0xb19d */
            {8'h00}, /* 0xb19c */
            {8'h00}, /* 0xb19b */
            {8'h00}, /* 0xb19a */
            {8'h00}, /* 0xb199 */
            {8'h00}, /* 0xb198 */
            {8'h00}, /* 0xb197 */
            {8'h00}, /* 0xb196 */
            {8'h00}, /* 0xb195 */
            {8'h00}, /* 0xb194 */
            {8'h00}, /* 0xb193 */
            {8'h00}, /* 0xb192 */
            {8'h00}, /* 0xb191 */
            {8'h00}, /* 0xb190 */
            {8'h00}, /* 0xb18f */
            {8'h00}, /* 0xb18e */
            {8'h00}, /* 0xb18d */
            {8'h00}, /* 0xb18c */
            {8'h00}, /* 0xb18b */
            {8'h00}, /* 0xb18a */
            {8'h00}, /* 0xb189 */
            {8'h00}, /* 0xb188 */
            {8'h00}, /* 0xb187 */
            {8'h00}, /* 0xb186 */
            {8'h00}, /* 0xb185 */
            {8'h00}, /* 0xb184 */
            {8'h00}, /* 0xb183 */
            {8'h00}, /* 0xb182 */
            {8'h00}, /* 0xb181 */
            {8'h00}, /* 0xb180 */
            {8'h00}, /* 0xb17f */
            {8'h00}, /* 0xb17e */
            {8'h00}, /* 0xb17d */
            {8'h00}, /* 0xb17c */
            {8'h00}, /* 0xb17b */
            {8'h00}, /* 0xb17a */
            {8'h00}, /* 0xb179 */
            {8'h00}, /* 0xb178 */
            {8'h00}, /* 0xb177 */
            {8'h00}, /* 0xb176 */
            {8'h00}, /* 0xb175 */
            {8'h00}, /* 0xb174 */
            {8'h00}, /* 0xb173 */
            {8'h00}, /* 0xb172 */
            {8'h00}, /* 0xb171 */
            {8'h00}, /* 0xb170 */
            {8'h00}, /* 0xb16f */
            {8'h00}, /* 0xb16e */
            {8'h00}, /* 0xb16d */
            {8'h00}, /* 0xb16c */
            {8'h00}, /* 0xb16b */
            {8'h00}, /* 0xb16a */
            {8'h00}, /* 0xb169 */
            {8'h00}, /* 0xb168 */
            {8'h00}, /* 0xb167 */
            {8'h00}, /* 0xb166 */
            {8'h00}, /* 0xb165 */
            {8'h00}, /* 0xb164 */
            {8'h00}, /* 0xb163 */
            {8'h00}, /* 0xb162 */
            {8'h00}, /* 0xb161 */
            {8'h00}, /* 0xb160 */
            {8'h00}, /* 0xb15f */
            {8'h00}, /* 0xb15e */
            {8'h00}, /* 0xb15d */
            {8'h00}, /* 0xb15c */
            {8'h00}, /* 0xb15b */
            {8'h00}, /* 0xb15a */
            {8'h00}, /* 0xb159 */
            {8'h00}, /* 0xb158 */
            {8'h00}, /* 0xb157 */
            {8'h00}, /* 0xb156 */
            {8'h00}, /* 0xb155 */
            {8'h00}, /* 0xb154 */
            {8'h00}, /* 0xb153 */
            {8'h00}, /* 0xb152 */
            {8'h00}, /* 0xb151 */
            {8'h00}, /* 0xb150 */
            {8'h00}, /* 0xb14f */
            {8'h00}, /* 0xb14e */
            {8'h00}, /* 0xb14d */
            {8'h00}, /* 0xb14c */
            {8'h00}, /* 0xb14b */
            {8'h00}, /* 0xb14a */
            {8'h00}, /* 0xb149 */
            {8'h00}, /* 0xb148 */
            {8'h00}, /* 0xb147 */
            {8'h00}, /* 0xb146 */
            {8'h00}, /* 0xb145 */
            {8'h00}, /* 0xb144 */
            {8'h00}, /* 0xb143 */
            {8'h00}, /* 0xb142 */
            {8'h00}, /* 0xb141 */
            {8'h00}, /* 0xb140 */
            {8'h00}, /* 0xb13f */
            {8'h00}, /* 0xb13e */
            {8'h00}, /* 0xb13d */
            {8'h00}, /* 0xb13c */
            {8'h00}, /* 0xb13b */
            {8'h00}, /* 0xb13a */
            {8'h00}, /* 0xb139 */
            {8'h00}, /* 0xb138 */
            {8'h00}, /* 0xb137 */
            {8'h00}, /* 0xb136 */
            {8'h00}, /* 0xb135 */
            {8'h00}, /* 0xb134 */
            {8'h00}, /* 0xb133 */
            {8'h00}, /* 0xb132 */
            {8'h00}, /* 0xb131 */
            {8'h00}, /* 0xb130 */
            {8'h00}, /* 0xb12f */
            {8'h00}, /* 0xb12e */
            {8'h00}, /* 0xb12d */
            {8'h00}, /* 0xb12c */
            {8'h00}, /* 0xb12b */
            {8'h00}, /* 0xb12a */
            {8'h00}, /* 0xb129 */
            {8'h00}, /* 0xb128 */
            {8'h00}, /* 0xb127 */
            {8'h00}, /* 0xb126 */
            {8'h00}, /* 0xb125 */
            {8'h00}, /* 0xb124 */
            {8'h00}, /* 0xb123 */
            {8'h00}, /* 0xb122 */
            {8'h00}, /* 0xb121 */
            {8'h00}, /* 0xb120 */
            {8'h00}, /* 0xb11f */
            {8'h00}, /* 0xb11e */
            {8'h00}, /* 0xb11d */
            {8'h00}, /* 0xb11c */
            {8'h00}, /* 0xb11b */
            {8'h00}, /* 0xb11a */
            {8'h00}, /* 0xb119 */
            {8'h00}, /* 0xb118 */
            {8'h00}, /* 0xb117 */
            {8'h00}, /* 0xb116 */
            {8'h00}, /* 0xb115 */
            {8'h00}, /* 0xb114 */
            {8'h00}, /* 0xb113 */
            {8'h00}, /* 0xb112 */
            {8'h00}, /* 0xb111 */
            {8'h00}, /* 0xb110 */
            {8'h00}, /* 0xb10f */
            {8'h00}, /* 0xb10e */
            {8'h00}, /* 0xb10d */
            {8'h00}, /* 0xb10c */
            {8'h00}, /* 0xb10b */
            {8'h00}, /* 0xb10a */
            {8'h00}, /* 0xb109 */
            {8'h00}, /* 0xb108 */
            {8'h00}, /* 0xb107 */
            {8'h00}, /* 0xb106 */
            {8'h00}, /* 0xb105 */
            {8'h00}, /* 0xb104 */
            {8'h00}, /* 0xb103 */
            {8'h00}, /* 0xb102 */
            {8'h00}, /* 0xb101 */
            {8'h00}, /* 0xb100 */
            {8'h00}, /* 0xb0ff */
            {8'h00}, /* 0xb0fe */
            {8'h00}, /* 0xb0fd */
            {8'h00}, /* 0xb0fc */
            {8'h00}, /* 0xb0fb */
            {8'h00}, /* 0xb0fa */
            {8'h00}, /* 0xb0f9 */
            {8'h00}, /* 0xb0f8 */
            {8'h00}, /* 0xb0f7 */
            {8'h00}, /* 0xb0f6 */
            {8'h00}, /* 0xb0f5 */
            {8'h00}, /* 0xb0f4 */
            {8'h00}, /* 0xb0f3 */
            {8'h00}, /* 0xb0f2 */
            {8'h00}, /* 0xb0f1 */
            {8'h00}, /* 0xb0f0 */
            {8'h00}, /* 0xb0ef */
            {8'h00}, /* 0xb0ee */
            {8'h00}, /* 0xb0ed */
            {8'h00}, /* 0xb0ec */
            {8'h00}, /* 0xb0eb */
            {8'h00}, /* 0xb0ea */
            {8'h00}, /* 0xb0e9 */
            {8'h00}, /* 0xb0e8 */
            {8'h00}, /* 0xb0e7 */
            {8'h00}, /* 0xb0e6 */
            {8'h00}, /* 0xb0e5 */
            {8'h00}, /* 0xb0e4 */
            {8'h00}, /* 0xb0e3 */
            {8'h00}, /* 0xb0e2 */
            {8'h00}, /* 0xb0e1 */
            {8'h00}, /* 0xb0e0 */
            {8'h00}, /* 0xb0df */
            {8'h00}, /* 0xb0de */
            {8'h00}, /* 0xb0dd */
            {8'h00}, /* 0xb0dc */
            {8'h00}, /* 0xb0db */
            {8'h00}, /* 0xb0da */
            {8'h00}, /* 0xb0d9 */
            {8'h00}, /* 0xb0d8 */
            {8'h00}, /* 0xb0d7 */
            {8'h00}, /* 0xb0d6 */
            {8'h00}, /* 0xb0d5 */
            {8'h00}, /* 0xb0d4 */
            {8'h00}, /* 0xb0d3 */
            {8'h00}, /* 0xb0d2 */
            {8'h00}, /* 0xb0d1 */
            {8'h00}, /* 0xb0d0 */
            {8'h00}, /* 0xb0cf */
            {8'h00}, /* 0xb0ce */
            {8'h00}, /* 0xb0cd */
            {8'h00}, /* 0xb0cc */
            {8'h00}, /* 0xb0cb */
            {8'h00}, /* 0xb0ca */
            {8'h00}, /* 0xb0c9 */
            {8'h00}, /* 0xb0c8 */
            {8'h00}, /* 0xb0c7 */
            {8'h00}, /* 0xb0c6 */
            {8'h00}, /* 0xb0c5 */
            {8'h00}, /* 0xb0c4 */
            {8'h00}, /* 0xb0c3 */
            {8'h00}, /* 0xb0c2 */
            {8'h00}, /* 0xb0c1 */
            {8'h00}, /* 0xb0c0 */
            {8'h00}, /* 0xb0bf */
            {8'h00}, /* 0xb0be */
            {8'h00}, /* 0xb0bd */
            {8'h00}, /* 0xb0bc */
            {8'h00}, /* 0xb0bb */
            {8'h00}, /* 0xb0ba */
            {8'h00}, /* 0xb0b9 */
            {8'h00}, /* 0xb0b8 */
            {8'h00}, /* 0xb0b7 */
            {8'h00}, /* 0xb0b6 */
            {8'h00}, /* 0xb0b5 */
            {8'h00}, /* 0xb0b4 */
            {8'h00}, /* 0xb0b3 */
            {8'h00}, /* 0xb0b2 */
            {8'h00}, /* 0xb0b1 */
            {8'h00}, /* 0xb0b0 */
            {8'h00}, /* 0xb0af */
            {8'h00}, /* 0xb0ae */
            {8'h00}, /* 0xb0ad */
            {8'h00}, /* 0xb0ac */
            {8'h00}, /* 0xb0ab */
            {8'h00}, /* 0xb0aa */
            {8'h00}, /* 0xb0a9 */
            {8'h00}, /* 0xb0a8 */
            {8'h00}, /* 0xb0a7 */
            {8'h00}, /* 0xb0a6 */
            {8'h00}, /* 0xb0a5 */
            {8'h00}, /* 0xb0a4 */
            {8'h00}, /* 0xb0a3 */
            {8'h00}, /* 0xb0a2 */
            {8'h00}, /* 0xb0a1 */
            {8'h00}, /* 0xb0a0 */
            {8'h00}, /* 0xb09f */
            {8'h00}, /* 0xb09e */
            {8'h00}, /* 0xb09d */
            {8'h00}, /* 0xb09c */
            {8'h00}, /* 0xb09b */
            {8'h00}, /* 0xb09a */
            {8'h00}, /* 0xb099 */
            {8'h00}, /* 0xb098 */
            {8'h00}, /* 0xb097 */
            {8'h00}, /* 0xb096 */
            {8'h00}, /* 0xb095 */
            {8'h00}, /* 0xb094 */
            {8'h00}, /* 0xb093 */
            {8'h00}, /* 0xb092 */
            {8'h00}, /* 0xb091 */
            {8'h00}, /* 0xb090 */
            {8'h00}, /* 0xb08f */
            {8'h00}, /* 0xb08e */
            {8'h00}, /* 0xb08d */
            {8'h00}, /* 0xb08c */
            {8'h00}, /* 0xb08b */
            {8'h00}, /* 0xb08a */
            {8'h00}, /* 0xb089 */
            {8'h00}, /* 0xb088 */
            {8'h00}, /* 0xb087 */
            {8'h00}, /* 0xb086 */
            {8'h00}, /* 0xb085 */
            {8'h00}, /* 0xb084 */
            {8'h00}, /* 0xb083 */
            {8'h00}, /* 0xb082 */
            {8'h00}, /* 0xb081 */
            {8'h00}, /* 0xb080 */
            {8'h00}, /* 0xb07f */
            {8'h00}, /* 0xb07e */
            {8'h00}, /* 0xb07d */
            {8'h00}, /* 0xb07c */
            {8'h00}, /* 0xb07b */
            {8'h00}, /* 0xb07a */
            {8'h00}, /* 0xb079 */
            {8'h00}, /* 0xb078 */
            {8'h00}, /* 0xb077 */
            {8'h00}, /* 0xb076 */
            {8'h00}, /* 0xb075 */
            {8'h00}, /* 0xb074 */
            {8'h00}, /* 0xb073 */
            {8'h00}, /* 0xb072 */
            {8'h00}, /* 0xb071 */
            {8'h00}, /* 0xb070 */
            {8'h00}, /* 0xb06f */
            {8'h00}, /* 0xb06e */
            {8'h00}, /* 0xb06d */
            {8'h00}, /* 0xb06c */
            {8'h00}, /* 0xb06b */
            {8'h00}, /* 0xb06a */
            {8'h00}, /* 0xb069 */
            {8'h00}, /* 0xb068 */
            {8'h00}, /* 0xb067 */
            {8'h00}, /* 0xb066 */
            {8'h00}, /* 0xb065 */
            {8'h00}, /* 0xb064 */
            {8'h00}, /* 0xb063 */
            {8'h00}, /* 0xb062 */
            {8'h00}, /* 0xb061 */
            {8'h00}, /* 0xb060 */
            {8'h00}, /* 0xb05f */
            {8'h00}, /* 0xb05e */
            {8'h00}, /* 0xb05d */
            {8'h00}, /* 0xb05c */
            {8'h00}, /* 0xb05b */
            {8'h00}, /* 0xb05a */
            {8'h00}, /* 0xb059 */
            {8'h00}, /* 0xb058 */
            {8'h00}, /* 0xb057 */
            {8'h00}, /* 0xb056 */
            {8'h00}, /* 0xb055 */
            {8'h00}, /* 0xb054 */
            {8'h00}, /* 0xb053 */
            {8'h00}, /* 0xb052 */
            {8'h00}, /* 0xb051 */
            {8'h00}, /* 0xb050 */
            {8'h00}, /* 0xb04f */
            {8'h00}, /* 0xb04e */
            {8'h00}, /* 0xb04d */
            {8'h00}, /* 0xb04c */
            {8'h00}, /* 0xb04b */
            {8'h00}, /* 0xb04a */
            {8'h00}, /* 0xb049 */
            {8'h00}, /* 0xb048 */
            {8'h00}, /* 0xb047 */
            {8'h00}, /* 0xb046 */
            {8'h00}, /* 0xb045 */
            {8'h00}, /* 0xb044 */
            {8'h00}, /* 0xb043 */
            {8'h00}, /* 0xb042 */
            {8'h00}, /* 0xb041 */
            {8'h00}, /* 0xb040 */
            {8'h00}, /* 0xb03f */
            {8'h00}, /* 0xb03e */
            {8'h00}, /* 0xb03d */
            {8'h00}, /* 0xb03c */
            {8'h00}, /* 0xb03b */
            {8'h00}, /* 0xb03a */
            {8'h00}, /* 0xb039 */
            {8'h00}, /* 0xb038 */
            {8'h00}, /* 0xb037 */
            {8'h00}, /* 0xb036 */
            {8'h00}, /* 0xb035 */
            {8'h00}, /* 0xb034 */
            {8'h00}, /* 0xb033 */
            {8'h00}, /* 0xb032 */
            {8'h00}, /* 0xb031 */
            {8'h00}, /* 0xb030 */
            {8'h00}, /* 0xb02f */
            {8'h00}, /* 0xb02e */
            {8'h00}, /* 0xb02d */
            {8'h00}, /* 0xb02c */
            {8'h00}, /* 0xb02b */
            {8'h00}, /* 0xb02a */
            {8'h00}, /* 0xb029 */
            {8'h00}, /* 0xb028 */
            {8'h00}, /* 0xb027 */
            {8'h00}, /* 0xb026 */
            {8'h00}, /* 0xb025 */
            {8'h00}, /* 0xb024 */
            {8'h00}, /* 0xb023 */
            {8'h00}, /* 0xb022 */
            {8'h00}, /* 0xb021 */
            {8'h00}, /* 0xb020 */
            {8'h00}, /* 0xb01f */
            {8'h00}, /* 0xb01e */
            {8'h00}, /* 0xb01d */
            {8'h00}, /* 0xb01c */
            {8'h00}, /* 0xb01b */
            {8'h00}, /* 0xb01a */
            {8'h00}, /* 0xb019 */
            {8'h00}, /* 0xb018 */
            {8'h00}, /* 0xb017 */
            {8'h00}, /* 0xb016 */
            {8'h00}, /* 0xb015 */
            {8'h00}, /* 0xb014 */
            {8'h00}, /* 0xb013 */
            {8'h00}, /* 0xb012 */
            {8'h00}, /* 0xb011 */
            {8'h00}, /* 0xb010 */
            {8'h00}, /* 0xb00f */
            {8'h00}, /* 0xb00e */
            {8'h00}, /* 0xb00d */
            {8'h00}, /* 0xb00c */
            {8'h00}, /* 0xb00b */
            {8'h00}, /* 0xb00a */
            {8'h00}, /* 0xb009 */
            {8'h00}, /* 0xb008 */
            {8'h00}, /* 0xb007 */
            {8'h00}, /* 0xb006 */
            {8'h00}, /* 0xb005 */
            {8'h00}, /* 0xb004 */
            {8'h00}, /* 0xb003 */
            {8'h00}, /* 0xb002 */
            {8'h00}, /* 0xb001 */
            {8'h00}, /* 0xb000 */
            {8'h00}, /* 0xafff */
            {8'h00}, /* 0xaffe */
            {8'h00}, /* 0xaffd */
            {8'h00}, /* 0xaffc */
            {8'h00}, /* 0xaffb */
            {8'h00}, /* 0xaffa */
            {8'h00}, /* 0xaff9 */
            {8'h00}, /* 0xaff8 */
            {8'h00}, /* 0xaff7 */
            {8'h00}, /* 0xaff6 */
            {8'h00}, /* 0xaff5 */
            {8'h00}, /* 0xaff4 */
            {8'h00}, /* 0xaff3 */
            {8'h00}, /* 0xaff2 */
            {8'h00}, /* 0xaff1 */
            {8'h00}, /* 0xaff0 */
            {8'h00}, /* 0xafef */
            {8'h00}, /* 0xafee */
            {8'h00}, /* 0xafed */
            {8'h00}, /* 0xafec */
            {8'h00}, /* 0xafeb */
            {8'h00}, /* 0xafea */
            {8'h00}, /* 0xafe9 */
            {8'h00}, /* 0xafe8 */
            {8'h00}, /* 0xafe7 */
            {8'h00}, /* 0xafe6 */
            {8'h00}, /* 0xafe5 */
            {8'h00}, /* 0xafe4 */
            {8'h00}, /* 0xafe3 */
            {8'h00}, /* 0xafe2 */
            {8'h00}, /* 0xafe1 */
            {8'h00}, /* 0xafe0 */
            {8'h00}, /* 0xafdf */
            {8'h00}, /* 0xafde */
            {8'h00}, /* 0xafdd */
            {8'h00}, /* 0xafdc */
            {8'h00}, /* 0xafdb */
            {8'h00}, /* 0xafda */
            {8'h00}, /* 0xafd9 */
            {8'h00}, /* 0xafd8 */
            {8'h00}, /* 0xafd7 */
            {8'h00}, /* 0xafd6 */
            {8'h00}, /* 0xafd5 */
            {8'h00}, /* 0xafd4 */
            {8'h00}, /* 0xafd3 */
            {8'h00}, /* 0xafd2 */
            {8'h00}, /* 0xafd1 */
            {8'h00}, /* 0xafd0 */
            {8'h00}, /* 0xafcf */
            {8'h00}, /* 0xafce */
            {8'h00}, /* 0xafcd */
            {8'h00}, /* 0xafcc */
            {8'h00}, /* 0xafcb */
            {8'h00}, /* 0xafca */
            {8'h00}, /* 0xafc9 */
            {8'h00}, /* 0xafc8 */
            {8'h00}, /* 0xafc7 */
            {8'h00}, /* 0xafc6 */
            {8'h00}, /* 0xafc5 */
            {8'h00}, /* 0xafc4 */
            {8'h00}, /* 0xafc3 */
            {8'h00}, /* 0xafc2 */
            {8'h00}, /* 0xafc1 */
            {8'h00}, /* 0xafc0 */
            {8'h00}, /* 0xafbf */
            {8'h00}, /* 0xafbe */
            {8'h00}, /* 0xafbd */
            {8'h00}, /* 0xafbc */
            {8'h00}, /* 0xafbb */
            {8'h00}, /* 0xafba */
            {8'h00}, /* 0xafb9 */
            {8'h00}, /* 0xafb8 */
            {8'h00}, /* 0xafb7 */
            {8'h00}, /* 0xafb6 */
            {8'h00}, /* 0xafb5 */
            {8'h00}, /* 0xafb4 */
            {8'h00}, /* 0xafb3 */
            {8'h00}, /* 0xafb2 */
            {8'h00}, /* 0xafb1 */
            {8'h00}, /* 0xafb0 */
            {8'h00}, /* 0xafaf */
            {8'h00}, /* 0xafae */
            {8'h00}, /* 0xafad */
            {8'h00}, /* 0xafac */
            {8'h00}, /* 0xafab */
            {8'h00}, /* 0xafaa */
            {8'h00}, /* 0xafa9 */
            {8'h00}, /* 0xafa8 */
            {8'h00}, /* 0xafa7 */
            {8'h00}, /* 0xafa6 */
            {8'h00}, /* 0xafa5 */
            {8'h00}, /* 0xafa4 */
            {8'h00}, /* 0xafa3 */
            {8'h00}, /* 0xafa2 */
            {8'h00}, /* 0xafa1 */
            {8'h00}, /* 0xafa0 */
            {8'h00}, /* 0xaf9f */
            {8'h00}, /* 0xaf9e */
            {8'h00}, /* 0xaf9d */
            {8'h00}, /* 0xaf9c */
            {8'h00}, /* 0xaf9b */
            {8'h00}, /* 0xaf9a */
            {8'h00}, /* 0xaf99 */
            {8'h00}, /* 0xaf98 */
            {8'h00}, /* 0xaf97 */
            {8'h00}, /* 0xaf96 */
            {8'h00}, /* 0xaf95 */
            {8'h00}, /* 0xaf94 */
            {8'h00}, /* 0xaf93 */
            {8'h00}, /* 0xaf92 */
            {8'h00}, /* 0xaf91 */
            {8'h00}, /* 0xaf90 */
            {8'h00}, /* 0xaf8f */
            {8'h00}, /* 0xaf8e */
            {8'h00}, /* 0xaf8d */
            {8'h00}, /* 0xaf8c */
            {8'h00}, /* 0xaf8b */
            {8'h00}, /* 0xaf8a */
            {8'h00}, /* 0xaf89 */
            {8'h00}, /* 0xaf88 */
            {8'h00}, /* 0xaf87 */
            {8'h00}, /* 0xaf86 */
            {8'h00}, /* 0xaf85 */
            {8'h00}, /* 0xaf84 */
            {8'h00}, /* 0xaf83 */
            {8'h00}, /* 0xaf82 */
            {8'h00}, /* 0xaf81 */
            {8'h00}, /* 0xaf80 */
            {8'h00}, /* 0xaf7f */
            {8'h00}, /* 0xaf7e */
            {8'h00}, /* 0xaf7d */
            {8'h00}, /* 0xaf7c */
            {8'h00}, /* 0xaf7b */
            {8'h00}, /* 0xaf7a */
            {8'h00}, /* 0xaf79 */
            {8'h00}, /* 0xaf78 */
            {8'h00}, /* 0xaf77 */
            {8'h00}, /* 0xaf76 */
            {8'h00}, /* 0xaf75 */
            {8'h00}, /* 0xaf74 */
            {8'h00}, /* 0xaf73 */
            {8'h00}, /* 0xaf72 */
            {8'h00}, /* 0xaf71 */
            {8'h00}, /* 0xaf70 */
            {8'h00}, /* 0xaf6f */
            {8'h00}, /* 0xaf6e */
            {8'h00}, /* 0xaf6d */
            {8'h00}, /* 0xaf6c */
            {8'h00}, /* 0xaf6b */
            {8'h00}, /* 0xaf6a */
            {8'h00}, /* 0xaf69 */
            {8'h00}, /* 0xaf68 */
            {8'h00}, /* 0xaf67 */
            {8'h00}, /* 0xaf66 */
            {8'h00}, /* 0xaf65 */
            {8'h00}, /* 0xaf64 */
            {8'h00}, /* 0xaf63 */
            {8'h00}, /* 0xaf62 */
            {8'h00}, /* 0xaf61 */
            {8'h00}, /* 0xaf60 */
            {8'h00}, /* 0xaf5f */
            {8'h00}, /* 0xaf5e */
            {8'h00}, /* 0xaf5d */
            {8'h00}, /* 0xaf5c */
            {8'h00}, /* 0xaf5b */
            {8'h00}, /* 0xaf5a */
            {8'h00}, /* 0xaf59 */
            {8'h00}, /* 0xaf58 */
            {8'h00}, /* 0xaf57 */
            {8'h00}, /* 0xaf56 */
            {8'h00}, /* 0xaf55 */
            {8'h00}, /* 0xaf54 */
            {8'h00}, /* 0xaf53 */
            {8'h00}, /* 0xaf52 */
            {8'h00}, /* 0xaf51 */
            {8'h00}, /* 0xaf50 */
            {8'h00}, /* 0xaf4f */
            {8'h00}, /* 0xaf4e */
            {8'h00}, /* 0xaf4d */
            {8'h00}, /* 0xaf4c */
            {8'h00}, /* 0xaf4b */
            {8'h00}, /* 0xaf4a */
            {8'h00}, /* 0xaf49 */
            {8'h00}, /* 0xaf48 */
            {8'h00}, /* 0xaf47 */
            {8'h00}, /* 0xaf46 */
            {8'h00}, /* 0xaf45 */
            {8'h00}, /* 0xaf44 */
            {8'h00}, /* 0xaf43 */
            {8'h00}, /* 0xaf42 */
            {8'h00}, /* 0xaf41 */
            {8'h00}, /* 0xaf40 */
            {8'h00}, /* 0xaf3f */
            {8'h00}, /* 0xaf3e */
            {8'h00}, /* 0xaf3d */
            {8'h00}, /* 0xaf3c */
            {8'h00}, /* 0xaf3b */
            {8'h00}, /* 0xaf3a */
            {8'h00}, /* 0xaf39 */
            {8'h00}, /* 0xaf38 */
            {8'h00}, /* 0xaf37 */
            {8'h00}, /* 0xaf36 */
            {8'h00}, /* 0xaf35 */
            {8'h00}, /* 0xaf34 */
            {8'h00}, /* 0xaf33 */
            {8'h00}, /* 0xaf32 */
            {8'h00}, /* 0xaf31 */
            {8'h00}, /* 0xaf30 */
            {8'h00}, /* 0xaf2f */
            {8'h00}, /* 0xaf2e */
            {8'h00}, /* 0xaf2d */
            {8'h00}, /* 0xaf2c */
            {8'h00}, /* 0xaf2b */
            {8'h00}, /* 0xaf2a */
            {8'h00}, /* 0xaf29 */
            {8'h00}, /* 0xaf28 */
            {8'h00}, /* 0xaf27 */
            {8'h00}, /* 0xaf26 */
            {8'h00}, /* 0xaf25 */
            {8'h00}, /* 0xaf24 */
            {8'h00}, /* 0xaf23 */
            {8'h00}, /* 0xaf22 */
            {8'h00}, /* 0xaf21 */
            {8'h00}, /* 0xaf20 */
            {8'h00}, /* 0xaf1f */
            {8'h00}, /* 0xaf1e */
            {8'h00}, /* 0xaf1d */
            {8'h00}, /* 0xaf1c */
            {8'h00}, /* 0xaf1b */
            {8'h00}, /* 0xaf1a */
            {8'h00}, /* 0xaf19 */
            {8'h00}, /* 0xaf18 */
            {8'h00}, /* 0xaf17 */
            {8'h00}, /* 0xaf16 */
            {8'h00}, /* 0xaf15 */
            {8'h00}, /* 0xaf14 */
            {8'h00}, /* 0xaf13 */
            {8'h00}, /* 0xaf12 */
            {8'h00}, /* 0xaf11 */
            {8'h00}, /* 0xaf10 */
            {8'h00}, /* 0xaf0f */
            {8'h00}, /* 0xaf0e */
            {8'h00}, /* 0xaf0d */
            {8'h00}, /* 0xaf0c */
            {8'h00}, /* 0xaf0b */
            {8'h00}, /* 0xaf0a */
            {8'h00}, /* 0xaf09 */
            {8'h00}, /* 0xaf08 */
            {8'h00}, /* 0xaf07 */
            {8'h00}, /* 0xaf06 */
            {8'h00}, /* 0xaf05 */
            {8'h00}, /* 0xaf04 */
            {8'h00}, /* 0xaf03 */
            {8'h00}, /* 0xaf02 */
            {8'h00}, /* 0xaf01 */
            {8'h00}, /* 0xaf00 */
            {8'h00}, /* 0xaeff */
            {8'h00}, /* 0xaefe */
            {8'h00}, /* 0xaefd */
            {8'h00}, /* 0xaefc */
            {8'h00}, /* 0xaefb */
            {8'h00}, /* 0xaefa */
            {8'h00}, /* 0xaef9 */
            {8'h00}, /* 0xaef8 */
            {8'h00}, /* 0xaef7 */
            {8'h00}, /* 0xaef6 */
            {8'h00}, /* 0xaef5 */
            {8'h00}, /* 0xaef4 */
            {8'h00}, /* 0xaef3 */
            {8'h00}, /* 0xaef2 */
            {8'h00}, /* 0xaef1 */
            {8'h00}, /* 0xaef0 */
            {8'h00}, /* 0xaeef */
            {8'h00}, /* 0xaeee */
            {8'h00}, /* 0xaeed */
            {8'h00}, /* 0xaeec */
            {8'h00}, /* 0xaeeb */
            {8'h00}, /* 0xaeea */
            {8'h00}, /* 0xaee9 */
            {8'h00}, /* 0xaee8 */
            {8'h00}, /* 0xaee7 */
            {8'h00}, /* 0xaee6 */
            {8'h00}, /* 0xaee5 */
            {8'h00}, /* 0xaee4 */
            {8'h00}, /* 0xaee3 */
            {8'h00}, /* 0xaee2 */
            {8'h00}, /* 0xaee1 */
            {8'h00}, /* 0xaee0 */
            {8'h00}, /* 0xaedf */
            {8'h00}, /* 0xaede */
            {8'h00}, /* 0xaedd */
            {8'h00}, /* 0xaedc */
            {8'h00}, /* 0xaedb */
            {8'h00}, /* 0xaeda */
            {8'h00}, /* 0xaed9 */
            {8'h00}, /* 0xaed8 */
            {8'h00}, /* 0xaed7 */
            {8'h00}, /* 0xaed6 */
            {8'h00}, /* 0xaed5 */
            {8'h00}, /* 0xaed4 */
            {8'h00}, /* 0xaed3 */
            {8'h00}, /* 0xaed2 */
            {8'h00}, /* 0xaed1 */
            {8'h00}, /* 0xaed0 */
            {8'h00}, /* 0xaecf */
            {8'h00}, /* 0xaece */
            {8'h00}, /* 0xaecd */
            {8'h00}, /* 0xaecc */
            {8'h00}, /* 0xaecb */
            {8'h00}, /* 0xaeca */
            {8'h00}, /* 0xaec9 */
            {8'h00}, /* 0xaec8 */
            {8'h00}, /* 0xaec7 */
            {8'h00}, /* 0xaec6 */
            {8'h00}, /* 0xaec5 */
            {8'h00}, /* 0xaec4 */
            {8'h00}, /* 0xaec3 */
            {8'h00}, /* 0xaec2 */
            {8'h00}, /* 0xaec1 */
            {8'h00}, /* 0xaec0 */
            {8'h00}, /* 0xaebf */
            {8'h00}, /* 0xaebe */
            {8'h00}, /* 0xaebd */
            {8'h00}, /* 0xaebc */
            {8'h00}, /* 0xaebb */
            {8'h00}, /* 0xaeba */
            {8'h00}, /* 0xaeb9 */
            {8'h00}, /* 0xaeb8 */
            {8'h00}, /* 0xaeb7 */
            {8'h00}, /* 0xaeb6 */
            {8'h00}, /* 0xaeb5 */
            {8'h00}, /* 0xaeb4 */
            {8'h00}, /* 0xaeb3 */
            {8'h00}, /* 0xaeb2 */
            {8'h00}, /* 0xaeb1 */
            {8'h00}, /* 0xaeb0 */
            {8'h00}, /* 0xaeaf */
            {8'h00}, /* 0xaeae */
            {8'h00}, /* 0xaead */
            {8'h00}, /* 0xaeac */
            {8'h00}, /* 0xaeab */
            {8'h00}, /* 0xaeaa */
            {8'h00}, /* 0xaea9 */
            {8'h00}, /* 0xaea8 */
            {8'h00}, /* 0xaea7 */
            {8'h00}, /* 0xaea6 */
            {8'h00}, /* 0xaea5 */
            {8'h00}, /* 0xaea4 */
            {8'h00}, /* 0xaea3 */
            {8'h00}, /* 0xaea2 */
            {8'h00}, /* 0xaea1 */
            {8'h00}, /* 0xaea0 */
            {8'h00}, /* 0xae9f */
            {8'h00}, /* 0xae9e */
            {8'h00}, /* 0xae9d */
            {8'h00}, /* 0xae9c */
            {8'h00}, /* 0xae9b */
            {8'h00}, /* 0xae9a */
            {8'h00}, /* 0xae99 */
            {8'h00}, /* 0xae98 */
            {8'h00}, /* 0xae97 */
            {8'h00}, /* 0xae96 */
            {8'h00}, /* 0xae95 */
            {8'h00}, /* 0xae94 */
            {8'h00}, /* 0xae93 */
            {8'h00}, /* 0xae92 */
            {8'h00}, /* 0xae91 */
            {8'h00}, /* 0xae90 */
            {8'h00}, /* 0xae8f */
            {8'h00}, /* 0xae8e */
            {8'h00}, /* 0xae8d */
            {8'h00}, /* 0xae8c */
            {8'h00}, /* 0xae8b */
            {8'h00}, /* 0xae8a */
            {8'h00}, /* 0xae89 */
            {8'h00}, /* 0xae88 */
            {8'h00}, /* 0xae87 */
            {8'h00}, /* 0xae86 */
            {8'h00}, /* 0xae85 */
            {8'h00}, /* 0xae84 */
            {8'h00}, /* 0xae83 */
            {8'h00}, /* 0xae82 */
            {8'h00}, /* 0xae81 */
            {8'h00}, /* 0xae80 */
            {8'h00}, /* 0xae7f */
            {8'h00}, /* 0xae7e */
            {8'h00}, /* 0xae7d */
            {8'h00}, /* 0xae7c */
            {8'h00}, /* 0xae7b */
            {8'h00}, /* 0xae7a */
            {8'h00}, /* 0xae79 */
            {8'h00}, /* 0xae78 */
            {8'h00}, /* 0xae77 */
            {8'h00}, /* 0xae76 */
            {8'h00}, /* 0xae75 */
            {8'h00}, /* 0xae74 */
            {8'h00}, /* 0xae73 */
            {8'h00}, /* 0xae72 */
            {8'h00}, /* 0xae71 */
            {8'h00}, /* 0xae70 */
            {8'h00}, /* 0xae6f */
            {8'h00}, /* 0xae6e */
            {8'h00}, /* 0xae6d */
            {8'h00}, /* 0xae6c */
            {8'h00}, /* 0xae6b */
            {8'h00}, /* 0xae6a */
            {8'h00}, /* 0xae69 */
            {8'h00}, /* 0xae68 */
            {8'h00}, /* 0xae67 */
            {8'h00}, /* 0xae66 */
            {8'h00}, /* 0xae65 */
            {8'h00}, /* 0xae64 */
            {8'h00}, /* 0xae63 */
            {8'h00}, /* 0xae62 */
            {8'h00}, /* 0xae61 */
            {8'h00}, /* 0xae60 */
            {8'h00}, /* 0xae5f */
            {8'h00}, /* 0xae5e */
            {8'h00}, /* 0xae5d */
            {8'h00}, /* 0xae5c */
            {8'h00}, /* 0xae5b */
            {8'h00}, /* 0xae5a */
            {8'h00}, /* 0xae59 */
            {8'h00}, /* 0xae58 */
            {8'h00}, /* 0xae57 */
            {8'h00}, /* 0xae56 */
            {8'h00}, /* 0xae55 */
            {8'h00}, /* 0xae54 */
            {8'h00}, /* 0xae53 */
            {8'h00}, /* 0xae52 */
            {8'h00}, /* 0xae51 */
            {8'h00}, /* 0xae50 */
            {8'h00}, /* 0xae4f */
            {8'h00}, /* 0xae4e */
            {8'h00}, /* 0xae4d */
            {8'h00}, /* 0xae4c */
            {8'h00}, /* 0xae4b */
            {8'h00}, /* 0xae4a */
            {8'h00}, /* 0xae49 */
            {8'h00}, /* 0xae48 */
            {8'h00}, /* 0xae47 */
            {8'h00}, /* 0xae46 */
            {8'h00}, /* 0xae45 */
            {8'h00}, /* 0xae44 */
            {8'h00}, /* 0xae43 */
            {8'h00}, /* 0xae42 */
            {8'h00}, /* 0xae41 */
            {8'h00}, /* 0xae40 */
            {8'h00}, /* 0xae3f */
            {8'h00}, /* 0xae3e */
            {8'h00}, /* 0xae3d */
            {8'h00}, /* 0xae3c */
            {8'h00}, /* 0xae3b */
            {8'h00}, /* 0xae3a */
            {8'h00}, /* 0xae39 */
            {8'h00}, /* 0xae38 */
            {8'h00}, /* 0xae37 */
            {8'h00}, /* 0xae36 */
            {8'h00}, /* 0xae35 */
            {8'h00}, /* 0xae34 */
            {8'h00}, /* 0xae33 */
            {8'h00}, /* 0xae32 */
            {8'h00}, /* 0xae31 */
            {8'h00}, /* 0xae30 */
            {8'h00}, /* 0xae2f */
            {8'h00}, /* 0xae2e */
            {8'h00}, /* 0xae2d */
            {8'h00}, /* 0xae2c */
            {8'h00}, /* 0xae2b */
            {8'h00}, /* 0xae2a */
            {8'h00}, /* 0xae29 */
            {8'h00}, /* 0xae28 */
            {8'h00}, /* 0xae27 */
            {8'h00}, /* 0xae26 */
            {8'h00}, /* 0xae25 */
            {8'h00}, /* 0xae24 */
            {8'h00}, /* 0xae23 */
            {8'h00}, /* 0xae22 */
            {8'h00}, /* 0xae21 */
            {8'h00}, /* 0xae20 */
            {8'h00}, /* 0xae1f */
            {8'h00}, /* 0xae1e */
            {8'h00}, /* 0xae1d */
            {8'h00}, /* 0xae1c */
            {8'h00}, /* 0xae1b */
            {8'h00}, /* 0xae1a */
            {8'h00}, /* 0xae19 */
            {8'h00}, /* 0xae18 */
            {8'h00}, /* 0xae17 */
            {8'h00}, /* 0xae16 */
            {8'h00}, /* 0xae15 */
            {8'h00}, /* 0xae14 */
            {8'h00}, /* 0xae13 */
            {8'h00}, /* 0xae12 */
            {8'h00}, /* 0xae11 */
            {8'h00}, /* 0xae10 */
            {8'h00}, /* 0xae0f */
            {8'h00}, /* 0xae0e */
            {8'h00}, /* 0xae0d */
            {8'h00}, /* 0xae0c */
            {8'h00}, /* 0xae0b */
            {8'h00}, /* 0xae0a */
            {8'h00}, /* 0xae09 */
            {8'h00}, /* 0xae08 */
            {8'h00}, /* 0xae07 */
            {8'h00}, /* 0xae06 */
            {8'h00}, /* 0xae05 */
            {8'h00}, /* 0xae04 */
            {8'h00}, /* 0xae03 */
            {8'h00}, /* 0xae02 */
            {8'h00}, /* 0xae01 */
            {8'h00}, /* 0xae00 */
            {8'h00}, /* 0xadff */
            {8'h00}, /* 0xadfe */
            {8'h00}, /* 0xadfd */
            {8'h00}, /* 0xadfc */
            {8'h00}, /* 0xadfb */
            {8'h00}, /* 0xadfa */
            {8'h00}, /* 0xadf9 */
            {8'h00}, /* 0xadf8 */
            {8'h00}, /* 0xadf7 */
            {8'h00}, /* 0xadf6 */
            {8'h00}, /* 0xadf5 */
            {8'h00}, /* 0xadf4 */
            {8'h00}, /* 0xadf3 */
            {8'h00}, /* 0xadf2 */
            {8'h00}, /* 0xadf1 */
            {8'h00}, /* 0xadf0 */
            {8'h00}, /* 0xadef */
            {8'h00}, /* 0xadee */
            {8'h00}, /* 0xaded */
            {8'h00}, /* 0xadec */
            {8'h00}, /* 0xadeb */
            {8'h00}, /* 0xadea */
            {8'h00}, /* 0xade9 */
            {8'h00}, /* 0xade8 */
            {8'h00}, /* 0xade7 */
            {8'h00}, /* 0xade6 */
            {8'h00}, /* 0xade5 */
            {8'h00}, /* 0xade4 */
            {8'h00}, /* 0xade3 */
            {8'h00}, /* 0xade2 */
            {8'h00}, /* 0xade1 */
            {8'h00}, /* 0xade0 */
            {8'h00}, /* 0xaddf */
            {8'h00}, /* 0xadde */
            {8'h00}, /* 0xaddd */
            {8'h00}, /* 0xaddc */
            {8'h00}, /* 0xaddb */
            {8'h00}, /* 0xadda */
            {8'h00}, /* 0xadd9 */
            {8'h00}, /* 0xadd8 */
            {8'h00}, /* 0xadd7 */
            {8'h00}, /* 0xadd6 */
            {8'h00}, /* 0xadd5 */
            {8'h00}, /* 0xadd4 */
            {8'h00}, /* 0xadd3 */
            {8'h00}, /* 0xadd2 */
            {8'h00}, /* 0xadd1 */
            {8'h00}, /* 0xadd0 */
            {8'h00}, /* 0xadcf */
            {8'h00}, /* 0xadce */
            {8'h00}, /* 0xadcd */
            {8'h00}, /* 0xadcc */
            {8'h00}, /* 0xadcb */
            {8'h00}, /* 0xadca */
            {8'h00}, /* 0xadc9 */
            {8'h00}, /* 0xadc8 */
            {8'h00}, /* 0xadc7 */
            {8'h00}, /* 0xadc6 */
            {8'h00}, /* 0xadc5 */
            {8'h00}, /* 0xadc4 */
            {8'h00}, /* 0xadc3 */
            {8'h00}, /* 0xadc2 */
            {8'h00}, /* 0xadc1 */
            {8'h00}, /* 0xadc0 */
            {8'h00}, /* 0xadbf */
            {8'h00}, /* 0xadbe */
            {8'h00}, /* 0xadbd */
            {8'h00}, /* 0xadbc */
            {8'h00}, /* 0xadbb */
            {8'h00}, /* 0xadba */
            {8'h00}, /* 0xadb9 */
            {8'h00}, /* 0xadb8 */
            {8'h00}, /* 0xadb7 */
            {8'h00}, /* 0xadb6 */
            {8'h00}, /* 0xadb5 */
            {8'h00}, /* 0xadb4 */
            {8'h00}, /* 0xadb3 */
            {8'h00}, /* 0xadb2 */
            {8'h00}, /* 0xadb1 */
            {8'h00}, /* 0xadb0 */
            {8'h00}, /* 0xadaf */
            {8'h00}, /* 0xadae */
            {8'h00}, /* 0xadad */
            {8'h00}, /* 0xadac */
            {8'h00}, /* 0xadab */
            {8'h00}, /* 0xadaa */
            {8'h00}, /* 0xada9 */
            {8'h00}, /* 0xada8 */
            {8'h00}, /* 0xada7 */
            {8'h00}, /* 0xada6 */
            {8'h00}, /* 0xada5 */
            {8'h00}, /* 0xada4 */
            {8'h00}, /* 0xada3 */
            {8'h00}, /* 0xada2 */
            {8'h00}, /* 0xada1 */
            {8'h00}, /* 0xada0 */
            {8'h00}, /* 0xad9f */
            {8'h00}, /* 0xad9e */
            {8'h00}, /* 0xad9d */
            {8'h00}, /* 0xad9c */
            {8'h00}, /* 0xad9b */
            {8'h00}, /* 0xad9a */
            {8'h00}, /* 0xad99 */
            {8'h00}, /* 0xad98 */
            {8'h00}, /* 0xad97 */
            {8'h00}, /* 0xad96 */
            {8'h00}, /* 0xad95 */
            {8'h00}, /* 0xad94 */
            {8'h00}, /* 0xad93 */
            {8'h00}, /* 0xad92 */
            {8'h00}, /* 0xad91 */
            {8'h00}, /* 0xad90 */
            {8'h00}, /* 0xad8f */
            {8'h00}, /* 0xad8e */
            {8'h00}, /* 0xad8d */
            {8'h00}, /* 0xad8c */
            {8'h00}, /* 0xad8b */
            {8'h00}, /* 0xad8a */
            {8'h00}, /* 0xad89 */
            {8'h00}, /* 0xad88 */
            {8'h00}, /* 0xad87 */
            {8'h00}, /* 0xad86 */
            {8'h00}, /* 0xad85 */
            {8'h00}, /* 0xad84 */
            {8'h00}, /* 0xad83 */
            {8'h00}, /* 0xad82 */
            {8'h00}, /* 0xad81 */
            {8'h00}, /* 0xad80 */
            {8'h00}, /* 0xad7f */
            {8'h00}, /* 0xad7e */
            {8'h00}, /* 0xad7d */
            {8'h00}, /* 0xad7c */
            {8'h00}, /* 0xad7b */
            {8'h00}, /* 0xad7a */
            {8'h00}, /* 0xad79 */
            {8'h00}, /* 0xad78 */
            {8'h00}, /* 0xad77 */
            {8'h00}, /* 0xad76 */
            {8'h00}, /* 0xad75 */
            {8'h00}, /* 0xad74 */
            {8'h00}, /* 0xad73 */
            {8'h00}, /* 0xad72 */
            {8'h00}, /* 0xad71 */
            {8'h00}, /* 0xad70 */
            {8'h00}, /* 0xad6f */
            {8'h00}, /* 0xad6e */
            {8'h00}, /* 0xad6d */
            {8'h00}, /* 0xad6c */
            {8'h00}, /* 0xad6b */
            {8'h00}, /* 0xad6a */
            {8'h00}, /* 0xad69 */
            {8'h00}, /* 0xad68 */
            {8'h00}, /* 0xad67 */
            {8'h00}, /* 0xad66 */
            {8'h00}, /* 0xad65 */
            {8'h00}, /* 0xad64 */
            {8'h00}, /* 0xad63 */
            {8'h00}, /* 0xad62 */
            {8'h00}, /* 0xad61 */
            {8'h00}, /* 0xad60 */
            {8'h00}, /* 0xad5f */
            {8'h00}, /* 0xad5e */
            {8'h00}, /* 0xad5d */
            {8'h00}, /* 0xad5c */
            {8'h00}, /* 0xad5b */
            {8'h00}, /* 0xad5a */
            {8'h00}, /* 0xad59 */
            {8'h00}, /* 0xad58 */
            {8'h00}, /* 0xad57 */
            {8'h00}, /* 0xad56 */
            {8'h00}, /* 0xad55 */
            {8'h00}, /* 0xad54 */
            {8'h00}, /* 0xad53 */
            {8'h00}, /* 0xad52 */
            {8'h00}, /* 0xad51 */
            {8'h00}, /* 0xad50 */
            {8'h00}, /* 0xad4f */
            {8'h00}, /* 0xad4e */
            {8'h00}, /* 0xad4d */
            {8'h00}, /* 0xad4c */
            {8'h00}, /* 0xad4b */
            {8'h00}, /* 0xad4a */
            {8'h00}, /* 0xad49 */
            {8'h00}, /* 0xad48 */
            {8'h00}, /* 0xad47 */
            {8'h00}, /* 0xad46 */
            {8'h00}, /* 0xad45 */
            {8'h00}, /* 0xad44 */
            {8'h00}, /* 0xad43 */
            {8'h00}, /* 0xad42 */
            {8'h00}, /* 0xad41 */
            {8'h00}, /* 0xad40 */
            {8'h00}, /* 0xad3f */
            {8'h00}, /* 0xad3e */
            {8'h00}, /* 0xad3d */
            {8'h00}, /* 0xad3c */
            {8'h00}, /* 0xad3b */
            {8'h00}, /* 0xad3a */
            {8'h00}, /* 0xad39 */
            {8'h00}, /* 0xad38 */
            {8'h00}, /* 0xad37 */
            {8'h00}, /* 0xad36 */
            {8'h00}, /* 0xad35 */
            {8'h00}, /* 0xad34 */
            {8'h00}, /* 0xad33 */
            {8'h00}, /* 0xad32 */
            {8'h00}, /* 0xad31 */
            {8'h00}, /* 0xad30 */
            {8'h00}, /* 0xad2f */
            {8'h00}, /* 0xad2e */
            {8'h00}, /* 0xad2d */
            {8'h00}, /* 0xad2c */
            {8'h00}, /* 0xad2b */
            {8'h00}, /* 0xad2a */
            {8'h00}, /* 0xad29 */
            {8'h00}, /* 0xad28 */
            {8'h00}, /* 0xad27 */
            {8'h00}, /* 0xad26 */
            {8'h00}, /* 0xad25 */
            {8'h00}, /* 0xad24 */
            {8'h00}, /* 0xad23 */
            {8'h00}, /* 0xad22 */
            {8'h00}, /* 0xad21 */
            {8'h00}, /* 0xad20 */
            {8'h00}, /* 0xad1f */
            {8'h00}, /* 0xad1e */
            {8'h00}, /* 0xad1d */
            {8'h00}, /* 0xad1c */
            {8'h00}, /* 0xad1b */
            {8'h00}, /* 0xad1a */
            {8'h00}, /* 0xad19 */
            {8'h00}, /* 0xad18 */
            {8'h00}, /* 0xad17 */
            {8'h00}, /* 0xad16 */
            {8'h00}, /* 0xad15 */
            {8'h00}, /* 0xad14 */
            {8'h00}, /* 0xad13 */
            {8'h00}, /* 0xad12 */
            {8'h00}, /* 0xad11 */
            {8'h00}, /* 0xad10 */
            {8'h00}, /* 0xad0f */
            {8'h00}, /* 0xad0e */
            {8'h00}, /* 0xad0d */
            {8'h00}, /* 0xad0c */
            {8'h00}, /* 0xad0b */
            {8'h00}, /* 0xad0a */
            {8'h00}, /* 0xad09 */
            {8'h00}, /* 0xad08 */
            {8'h00}, /* 0xad07 */
            {8'h00}, /* 0xad06 */
            {8'h00}, /* 0xad05 */
            {8'h00}, /* 0xad04 */
            {8'h00}, /* 0xad03 */
            {8'h00}, /* 0xad02 */
            {8'h00}, /* 0xad01 */
            {8'h00}, /* 0xad00 */
            {8'h00}, /* 0xacff */
            {8'h00}, /* 0xacfe */
            {8'h00}, /* 0xacfd */
            {8'h00}, /* 0xacfc */
            {8'h00}, /* 0xacfb */
            {8'h00}, /* 0xacfa */
            {8'h00}, /* 0xacf9 */
            {8'h00}, /* 0xacf8 */
            {8'h00}, /* 0xacf7 */
            {8'h00}, /* 0xacf6 */
            {8'h00}, /* 0xacf5 */
            {8'h00}, /* 0xacf4 */
            {8'h00}, /* 0xacf3 */
            {8'h00}, /* 0xacf2 */
            {8'h00}, /* 0xacf1 */
            {8'h00}, /* 0xacf0 */
            {8'h00}, /* 0xacef */
            {8'h00}, /* 0xacee */
            {8'h00}, /* 0xaced */
            {8'h00}, /* 0xacec */
            {8'h00}, /* 0xaceb */
            {8'h00}, /* 0xacea */
            {8'h00}, /* 0xace9 */
            {8'h00}, /* 0xace8 */
            {8'h00}, /* 0xace7 */
            {8'h00}, /* 0xace6 */
            {8'h00}, /* 0xace5 */
            {8'h00}, /* 0xace4 */
            {8'h00}, /* 0xace3 */
            {8'h00}, /* 0xace2 */
            {8'h00}, /* 0xace1 */
            {8'h00}, /* 0xace0 */
            {8'h00}, /* 0xacdf */
            {8'h00}, /* 0xacde */
            {8'h00}, /* 0xacdd */
            {8'h00}, /* 0xacdc */
            {8'h00}, /* 0xacdb */
            {8'h00}, /* 0xacda */
            {8'h00}, /* 0xacd9 */
            {8'h00}, /* 0xacd8 */
            {8'h00}, /* 0xacd7 */
            {8'h00}, /* 0xacd6 */
            {8'h00}, /* 0xacd5 */
            {8'h00}, /* 0xacd4 */
            {8'h00}, /* 0xacd3 */
            {8'h00}, /* 0xacd2 */
            {8'h00}, /* 0xacd1 */
            {8'h00}, /* 0xacd0 */
            {8'h00}, /* 0xaccf */
            {8'h00}, /* 0xacce */
            {8'h00}, /* 0xaccd */
            {8'h00}, /* 0xaccc */
            {8'h00}, /* 0xaccb */
            {8'h00}, /* 0xacca */
            {8'h00}, /* 0xacc9 */
            {8'h00}, /* 0xacc8 */
            {8'h00}, /* 0xacc7 */
            {8'h00}, /* 0xacc6 */
            {8'h00}, /* 0xacc5 */
            {8'h00}, /* 0xacc4 */
            {8'h00}, /* 0xacc3 */
            {8'h00}, /* 0xacc2 */
            {8'h00}, /* 0xacc1 */
            {8'h00}, /* 0xacc0 */
            {8'h00}, /* 0xacbf */
            {8'h00}, /* 0xacbe */
            {8'h00}, /* 0xacbd */
            {8'h00}, /* 0xacbc */
            {8'h00}, /* 0xacbb */
            {8'h00}, /* 0xacba */
            {8'h00}, /* 0xacb9 */
            {8'h00}, /* 0xacb8 */
            {8'h00}, /* 0xacb7 */
            {8'h00}, /* 0xacb6 */
            {8'h00}, /* 0xacb5 */
            {8'h00}, /* 0xacb4 */
            {8'h00}, /* 0xacb3 */
            {8'h00}, /* 0xacb2 */
            {8'h00}, /* 0xacb1 */
            {8'h00}, /* 0xacb0 */
            {8'h00}, /* 0xacaf */
            {8'h00}, /* 0xacae */
            {8'h00}, /* 0xacad */
            {8'h00}, /* 0xacac */
            {8'h00}, /* 0xacab */
            {8'h00}, /* 0xacaa */
            {8'h00}, /* 0xaca9 */
            {8'h00}, /* 0xaca8 */
            {8'h00}, /* 0xaca7 */
            {8'h00}, /* 0xaca6 */
            {8'h00}, /* 0xaca5 */
            {8'h00}, /* 0xaca4 */
            {8'h00}, /* 0xaca3 */
            {8'h00}, /* 0xaca2 */
            {8'h00}, /* 0xaca1 */
            {8'h00}, /* 0xaca0 */
            {8'h00}, /* 0xac9f */
            {8'h00}, /* 0xac9e */
            {8'h00}, /* 0xac9d */
            {8'h00}, /* 0xac9c */
            {8'h00}, /* 0xac9b */
            {8'h00}, /* 0xac9a */
            {8'h00}, /* 0xac99 */
            {8'h00}, /* 0xac98 */
            {8'h00}, /* 0xac97 */
            {8'h00}, /* 0xac96 */
            {8'h00}, /* 0xac95 */
            {8'h00}, /* 0xac94 */
            {8'h00}, /* 0xac93 */
            {8'h00}, /* 0xac92 */
            {8'h00}, /* 0xac91 */
            {8'h00}, /* 0xac90 */
            {8'h00}, /* 0xac8f */
            {8'h00}, /* 0xac8e */
            {8'h00}, /* 0xac8d */
            {8'h00}, /* 0xac8c */
            {8'h00}, /* 0xac8b */
            {8'h00}, /* 0xac8a */
            {8'h00}, /* 0xac89 */
            {8'h00}, /* 0xac88 */
            {8'h00}, /* 0xac87 */
            {8'h00}, /* 0xac86 */
            {8'h00}, /* 0xac85 */
            {8'h00}, /* 0xac84 */
            {8'h00}, /* 0xac83 */
            {8'h00}, /* 0xac82 */
            {8'h00}, /* 0xac81 */
            {8'h00}, /* 0xac80 */
            {8'h00}, /* 0xac7f */
            {8'h00}, /* 0xac7e */
            {8'h00}, /* 0xac7d */
            {8'h00}, /* 0xac7c */
            {8'h00}, /* 0xac7b */
            {8'h00}, /* 0xac7a */
            {8'h00}, /* 0xac79 */
            {8'h00}, /* 0xac78 */
            {8'h00}, /* 0xac77 */
            {8'h00}, /* 0xac76 */
            {8'h00}, /* 0xac75 */
            {8'h00}, /* 0xac74 */
            {8'h00}, /* 0xac73 */
            {8'h00}, /* 0xac72 */
            {8'h00}, /* 0xac71 */
            {8'h00}, /* 0xac70 */
            {8'h00}, /* 0xac6f */
            {8'h00}, /* 0xac6e */
            {8'h00}, /* 0xac6d */
            {8'h00}, /* 0xac6c */
            {8'h00}, /* 0xac6b */
            {8'h00}, /* 0xac6a */
            {8'h00}, /* 0xac69 */
            {8'h00}, /* 0xac68 */
            {8'h00}, /* 0xac67 */
            {8'h00}, /* 0xac66 */
            {8'h00}, /* 0xac65 */
            {8'h00}, /* 0xac64 */
            {8'h00}, /* 0xac63 */
            {8'h00}, /* 0xac62 */
            {8'h00}, /* 0xac61 */
            {8'h00}, /* 0xac60 */
            {8'h00}, /* 0xac5f */
            {8'h00}, /* 0xac5e */
            {8'h00}, /* 0xac5d */
            {8'h00}, /* 0xac5c */
            {8'h00}, /* 0xac5b */
            {8'h00}, /* 0xac5a */
            {8'h00}, /* 0xac59 */
            {8'h00}, /* 0xac58 */
            {8'h00}, /* 0xac57 */
            {8'h00}, /* 0xac56 */
            {8'h00}, /* 0xac55 */
            {8'h00}, /* 0xac54 */
            {8'h00}, /* 0xac53 */
            {8'h00}, /* 0xac52 */
            {8'h00}, /* 0xac51 */
            {8'h00}, /* 0xac50 */
            {8'h00}, /* 0xac4f */
            {8'h00}, /* 0xac4e */
            {8'h00}, /* 0xac4d */
            {8'h00}, /* 0xac4c */
            {8'h00}, /* 0xac4b */
            {8'h00}, /* 0xac4a */
            {8'h00}, /* 0xac49 */
            {8'h00}, /* 0xac48 */
            {8'h00}, /* 0xac47 */
            {8'h00}, /* 0xac46 */
            {8'h00}, /* 0xac45 */
            {8'h00}, /* 0xac44 */
            {8'h00}, /* 0xac43 */
            {8'h00}, /* 0xac42 */
            {8'h00}, /* 0xac41 */
            {8'h00}, /* 0xac40 */
            {8'h00}, /* 0xac3f */
            {8'h00}, /* 0xac3e */
            {8'h00}, /* 0xac3d */
            {8'h00}, /* 0xac3c */
            {8'h00}, /* 0xac3b */
            {8'h00}, /* 0xac3a */
            {8'h00}, /* 0xac39 */
            {8'h00}, /* 0xac38 */
            {8'h00}, /* 0xac37 */
            {8'h00}, /* 0xac36 */
            {8'h00}, /* 0xac35 */
            {8'h00}, /* 0xac34 */
            {8'h00}, /* 0xac33 */
            {8'h00}, /* 0xac32 */
            {8'h00}, /* 0xac31 */
            {8'h00}, /* 0xac30 */
            {8'h00}, /* 0xac2f */
            {8'h00}, /* 0xac2e */
            {8'h00}, /* 0xac2d */
            {8'h00}, /* 0xac2c */
            {8'h00}, /* 0xac2b */
            {8'h00}, /* 0xac2a */
            {8'h00}, /* 0xac29 */
            {8'h00}, /* 0xac28 */
            {8'h00}, /* 0xac27 */
            {8'h00}, /* 0xac26 */
            {8'h00}, /* 0xac25 */
            {8'h00}, /* 0xac24 */
            {8'h00}, /* 0xac23 */
            {8'h00}, /* 0xac22 */
            {8'h00}, /* 0xac21 */
            {8'h00}, /* 0xac20 */
            {8'h00}, /* 0xac1f */
            {8'h00}, /* 0xac1e */
            {8'h00}, /* 0xac1d */
            {8'h00}, /* 0xac1c */
            {8'h00}, /* 0xac1b */
            {8'h00}, /* 0xac1a */
            {8'h00}, /* 0xac19 */
            {8'h00}, /* 0xac18 */
            {8'h00}, /* 0xac17 */
            {8'h00}, /* 0xac16 */
            {8'h00}, /* 0xac15 */
            {8'h00}, /* 0xac14 */
            {8'h00}, /* 0xac13 */
            {8'h00}, /* 0xac12 */
            {8'h00}, /* 0xac11 */
            {8'h00}, /* 0xac10 */
            {8'h00}, /* 0xac0f */
            {8'h00}, /* 0xac0e */
            {8'h00}, /* 0xac0d */
            {8'h00}, /* 0xac0c */
            {8'h00}, /* 0xac0b */
            {8'h00}, /* 0xac0a */
            {8'h00}, /* 0xac09 */
            {8'h00}, /* 0xac08 */
            {8'h00}, /* 0xac07 */
            {8'h00}, /* 0xac06 */
            {8'h00}, /* 0xac05 */
            {8'h00}, /* 0xac04 */
            {8'h00}, /* 0xac03 */
            {8'h00}, /* 0xac02 */
            {8'h00}, /* 0xac01 */
            {8'h00}, /* 0xac00 */
            {8'h00}, /* 0xabff */
            {8'h00}, /* 0xabfe */
            {8'h00}, /* 0xabfd */
            {8'h00}, /* 0xabfc */
            {8'h00}, /* 0xabfb */
            {8'h00}, /* 0xabfa */
            {8'h00}, /* 0xabf9 */
            {8'h00}, /* 0xabf8 */
            {8'h00}, /* 0xabf7 */
            {8'h00}, /* 0xabf6 */
            {8'h00}, /* 0xabf5 */
            {8'h00}, /* 0xabf4 */
            {8'h00}, /* 0xabf3 */
            {8'h00}, /* 0xabf2 */
            {8'h00}, /* 0xabf1 */
            {8'h00}, /* 0xabf0 */
            {8'h00}, /* 0xabef */
            {8'h00}, /* 0xabee */
            {8'h00}, /* 0xabed */
            {8'h00}, /* 0xabec */
            {8'h00}, /* 0xabeb */
            {8'h00}, /* 0xabea */
            {8'h00}, /* 0xabe9 */
            {8'h00}, /* 0xabe8 */
            {8'h00}, /* 0xabe7 */
            {8'h00}, /* 0xabe6 */
            {8'h00}, /* 0xabe5 */
            {8'h00}, /* 0xabe4 */
            {8'h00}, /* 0xabe3 */
            {8'h00}, /* 0xabe2 */
            {8'h00}, /* 0xabe1 */
            {8'h00}, /* 0xabe0 */
            {8'h00}, /* 0xabdf */
            {8'h00}, /* 0xabde */
            {8'h00}, /* 0xabdd */
            {8'h00}, /* 0xabdc */
            {8'h00}, /* 0xabdb */
            {8'h00}, /* 0xabda */
            {8'h00}, /* 0xabd9 */
            {8'h00}, /* 0xabd8 */
            {8'h00}, /* 0xabd7 */
            {8'h00}, /* 0xabd6 */
            {8'h00}, /* 0xabd5 */
            {8'h00}, /* 0xabd4 */
            {8'h00}, /* 0xabd3 */
            {8'h00}, /* 0xabd2 */
            {8'h00}, /* 0xabd1 */
            {8'h00}, /* 0xabd0 */
            {8'h00}, /* 0xabcf */
            {8'h00}, /* 0xabce */
            {8'h00}, /* 0xabcd */
            {8'h00}, /* 0xabcc */
            {8'h00}, /* 0xabcb */
            {8'h00}, /* 0xabca */
            {8'h00}, /* 0xabc9 */
            {8'h00}, /* 0xabc8 */
            {8'h00}, /* 0xabc7 */
            {8'h00}, /* 0xabc6 */
            {8'h00}, /* 0xabc5 */
            {8'h00}, /* 0xabc4 */
            {8'h00}, /* 0xabc3 */
            {8'h00}, /* 0xabc2 */
            {8'h00}, /* 0xabc1 */
            {8'h00}, /* 0xabc0 */
            {8'h00}, /* 0xabbf */
            {8'h00}, /* 0xabbe */
            {8'h00}, /* 0xabbd */
            {8'h00}, /* 0xabbc */
            {8'h00}, /* 0xabbb */
            {8'h00}, /* 0xabba */
            {8'h00}, /* 0xabb9 */
            {8'h00}, /* 0xabb8 */
            {8'h00}, /* 0xabb7 */
            {8'h00}, /* 0xabb6 */
            {8'h00}, /* 0xabb5 */
            {8'h00}, /* 0xabb4 */
            {8'h00}, /* 0xabb3 */
            {8'h00}, /* 0xabb2 */
            {8'h00}, /* 0xabb1 */
            {8'h00}, /* 0xabb0 */
            {8'h00}, /* 0xabaf */
            {8'h00}, /* 0xabae */
            {8'h00}, /* 0xabad */
            {8'h00}, /* 0xabac */
            {8'h00}, /* 0xabab */
            {8'h00}, /* 0xabaa */
            {8'h00}, /* 0xaba9 */
            {8'h00}, /* 0xaba8 */
            {8'h00}, /* 0xaba7 */
            {8'h00}, /* 0xaba6 */
            {8'h00}, /* 0xaba5 */
            {8'h00}, /* 0xaba4 */
            {8'h00}, /* 0xaba3 */
            {8'h00}, /* 0xaba2 */
            {8'h00}, /* 0xaba1 */
            {8'h00}, /* 0xaba0 */
            {8'h00}, /* 0xab9f */
            {8'h00}, /* 0xab9e */
            {8'h00}, /* 0xab9d */
            {8'h00}, /* 0xab9c */
            {8'h00}, /* 0xab9b */
            {8'h00}, /* 0xab9a */
            {8'h00}, /* 0xab99 */
            {8'h00}, /* 0xab98 */
            {8'h00}, /* 0xab97 */
            {8'h00}, /* 0xab96 */
            {8'h00}, /* 0xab95 */
            {8'h00}, /* 0xab94 */
            {8'h00}, /* 0xab93 */
            {8'h00}, /* 0xab92 */
            {8'h00}, /* 0xab91 */
            {8'h00}, /* 0xab90 */
            {8'h00}, /* 0xab8f */
            {8'h00}, /* 0xab8e */
            {8'h00}, /* 0xab8d */
            {8'h00}, /* 0xab8c */
            {8'h00}, /* 0xab8b */
            {8'h00}, /* 0xab8a */
            {8'h00}, /* 0xab89 */
            {8'h00}, /* 0xab88 */
            {8'h00}, /* 0xab87 */
            {8'h00}, /* 0xab86 */
            {8'h00}, /* 0xab85 */
            {8'h00}, /* 0xab84 */
            {8'h00}, /* 0xab83 */
            {8'h00}, /* 0xab82 */
            {8'h00}, /* 0xab81 */
            {8'h00}, /* 0xab80 */
            {8'h00}, /* 0xab7f */
            {8'h00}, /* 0xab7e */
            {8'h00}, /* 0xab7d */
            {8'h00}, /* 0xab7c */
            {8'h00}, /* 0xab7b */
            {8'h00}, /* 0xab7a */
            {8'h00}, /* 0xab79 */
            {8'h00}, /* 0xab78 */
            {8'h00}, /* 0xab77 */
            {8'h00}, /* 0xab76 */
            {8'h00}, /* 0xab75 */
            {8'h00}, /* 0xab74 */
            {8'h00}, /* 0xab73 */
            {8'h00}, /* 0xab72 */
            {8'h00}, /* 0xab71 */
            {8'h00}, /* 0xab70 */
            {8'h00}, /* 0xab6f */
            {8'h00}, /* 0xab6e */
            {8'h00}, /* 0xab6d */
            {8'h00}, /* 0xab6c */
            {8'h00}, /* 0xab6b */
            {8'h00}, /* 0xab6a */
            {8'h00}, /* 0xab69 */
            {8'h00}, /* 0xab68 */
            {8'h00}, /* 0xab67 */
            {8'h00}, /* 0xab66 */
            {8'h00}, /* 0xab65 */
            {8'h00}, /* 0xab64 */
            {8'h00}, /* 0xab63 */
            {8'h00}, /* 0xab62 */
            {8'h00}, /* 0xab61 */
            {8'h00}, /* 0xab60 */
            {8'h00}, /* 0xab5f */
            {8'h00}, /* 0xab5e */
            {8'h00}, /* 0xab5d */
            {8'h00}, /* 0xab5c */
            {8'h00}, /* 0xab5b */
            {8'h00}, /* 0xab5a */
            {8'h00}, /* 0xab59 */
            {8'h00}, /* 0xab58 */
            {8'h00}, /* 0xab57 */
            {8'h00}, /* 0xab56 */
            {8'h00}, /* 0xab55 */
            {8'h00}, /* 0xab54 */
            {8'h00}, /* 0xab53 */
            {8'h00}, /* 0xab52 */
            {8'h00}, /* 0xab51 */
            {8'h00}, /* 0xab50 */
            {8'h00}, /* 0xab4f */
            {8'h00}, /* 0xab4e */
            {8'h00}, /* 0xab4d */
            {8'h00}, /* 0xab4c */
            {8'h00}, /* 0xab4b */
            {8'h00}, /* 0xab4a */
            {8'h00}, /* 0xab49 */
            {8'h00}, /* 0xab48 */
            {8'h00}, /* 0xab47 */
            {8'h00}, /* 0xab46 */
            {8'h00}, /* 0xab45 */
            {8'h00}, /* 0xab44 */
            {8'h00}, /* 0xab43 */
            {8'h00}, /* 0xab42 */
            {8'h00}, /* 0xab41 */
            {8'h00}, /* 0xab40 */
            {8'h00}, /* 0xab3f */
            {8'h00}, /* 0xab3e */
            {8'h00}, /* 0xab3d */
            {8'h00}, /* 0xab3c */
            {8'h00}, /* 0xab3b */
            {8'h00}, /* 0xab3a */
            {8'h00}, /* 0xab39 */
            {8'h00}, /* 0xab38 */
            {8'h00}, /* 0xab37 */
            {8'h00}, /* 0xab36 */
            {8'h00}, /* 0xab35 */
            {8'h00}, /* 0xab34 */
            {8'h00}, /* 0xab33 */
            {8'h00}, /* 0xab32 */
            {8'h00}, /* 0xab31 */
            {8'h00}, /* 0xab30 */
            {8'h00}, /* 0xab2f */
            {8'h00}, /* 0xab2e */
            {8'h00}, /* 0xab2d */
            {8'h00}, /* 0xab2c */
            {8'h00}, /* 0xab2b */
            {8'h00}, /* 0xab2a */
            {8'h00}, /* 0xab29 */
            {8'h00}, /* 0xab28 */
            {8'h00}, /* 0xab27 */
            {8'h00}, /* 0xab26 */
            {8'h00}, /* 0xab25 */
            {8'h00}, /* 0xab24 */
            {8'h00}, /* 0xab23 */
            {8'h00}, /* 0xab22 */
            {8'h00}, /* 0xab21 */
            {8'h00}, /* 0xab20 */
            {8'h00}, /* 0xab1f */
            {8'h00}, /* 0xab1e */
            {8'h00}, /* 0xab1d */
            {8'h00}, /* 0xab1c */
            {8'h00}, /* 0xab1b */
            {8'h00}, /* 0xab1a */
            {8'h00}, /* 0xab19 */
            {8'h00}, /* 0xab18 */
            {8'h00}, /* 0xab17 */
            {8'h00}, /* 0xab16 */
            {8'h00}, /* 0xab15 */
            {8'h00}, /* 0xab14 */
            {8'h00}, /* 0xab13 */
            {8'h00}, /* 0xab12 */
            {8'h00}, /* 0xab11 */
            {8'h00}, /* 0xab10 */
            {8'h00}, /* 0xab0f */
            {8'h00}, /* 0xab0e */
            {8'h00}, /* 0xab0d */
            {8'h00}, /* 0xab0c */
            {8'h00}, /* 0xab0b */
            {8'h00}, /* 0xab0a */
            {8'h00}, /* 0xab09 */
            {8'h00}, /* 0xab08 */
            {8'h00}, /* 0xab07 */
            {8'h00}, /* 0xab06 */
            {8'h00}, /* 0xab05 */
            {8'h00}, /* 0xab04 */
            {8'h00}, /* 0xab03 */
            {8'h00}, /* 0xab02 */
            {8'h00}, /* 0xab01 */
            {8'h00}, /* 0xab00 */
            {8'h00}, /* 0xaaff */
            {8'h00}, /* 0xaafe */
            {8'h00}, /* 0xaafd */
            {8'h00}, /* 0xaafc */
            {8'h00}, /* 0xaafb */
            {8'h00}, /* 0xaafa */
            {8'h00}, /* 0xaaf9 */
            {8'h00}, /* 0xaaf8 */
            {8'h00}, /* 0xaaf7 */
            {8'h00}, /* 0xaaf6 */
            {8'h00}, /* 0xaaf5 */
            {8'h00}, /* 0xaaf4 */
            {8'h00}, /* 0xaaf3 */
            {8'h00}, /* 0xaaf2 */
            {8'h00}, /* 0xaaf1 */
            {8'h00}, /* 0xaaf0 */
            {8'h00}, /* 0xaaef */
            {8'h00}, /* 0xaaee */
            {8'h00}, /* 0xaaed */
            {8'h00}, /* 0xaaec */
            {8'h00}, /* 0xaaeb */
            {8'h00}, /* 0xaaea */
            {8'h00}, /* 0xaae9 */
            {8'h00}, /* 0xaae8 */
            {8'h00}, /* 0xaae7 */
            {8'h00}, /* 0xaae6 */
            {8'h00}, /* 0xaae5 */
            {8'h00}, /* 0xaae4 */
            {8'h00}, /* 0xaae3 */
            {8'h00}, /* 0xaae2 */
            {8'h00}, /* 0xaae1 */
            {8'h00}, /* 0xaae0 */
            {8'h00}, /* 0xaadf */
            {8'h00}, /* 0xaade */
            {8'h00}, /* 0xaadd */
            {8'h00}, /* 0xaadc */
            {8'h00}, /* 0xaadb */
            {8'h00}, /* 0xaada */
            {8'h00}, /* 0xaad9 */
            {8'h00}, /* 0xaad8 */
            {8'h00}, /* 0xaad7 */
            {8'h00}, /* 0xaad6 */
            {8'h00}, /* 0xaad5 */
            {8'h00}, /* 0xaad4 */
            {8'h00}, /* 0xaad3 */
            {8'h00}, /* 0xaad2 */
            {8'h00}, /* 0xaad1 */
            {8'h00}, /* 0xaad0 */
            {8'h00}, /* 0xaacf */
            {8'h00}, /* 0xaace */
            {8'h00}, /* 0xaacd */
            {8'h00}, /* 0xaacc */
            {8'h00}, /* 0xaacb */
            {8'h00}, /* 0xaaca */
            {8'h00}, /* 0xaac9 */
            {8'h00}, /* 0xaac8 */
            {8'h00}, /* 0xaac7 */
            {8'h00}, /* 0xaac6 */
            {8'h00}, /* 0xaac5 */
            {8'h00}, /* 0xaac4 */
            {8'h00}, /* 0xaac3 */
            {8'h00}, /* 0xaac2 */
            {8'h00}, /* 0xaac1 */
            {8'h00}, /* 0xaac0 */
            {8'h00}, /* 0xaabf */
            {8'h00}, /* 0xaabe */
            {8'h00}, /* 0xaabd */
            {8'h00}, /* 0xaabc */
            {8'h00}, /* 0xaabb */
            {8'h00}, /* 0xaaba */
            {8'h00}, /* 0xaab9 */
            {8'h00}, /* 0xaab8 */
            {8'h00}, /* 0xaab7 */
            {8'h00}, /* 0xaab6 */
            {8'h00}, /* 0xaab5 */
            {8'h00}, /* 0xaab4 */
            {8'h00}, /* 0xaab3 */
            {8'h00}, /* 0xaab2 */
            {8'h00}, /* 0xaab1 */
            {8'h00}, /* 0xaab0 */
            {8'h00}, /* 0xaaaf */
            {8'h00}, /* 0xaaae */
            {8'h00}, /* 0xaaad */
            {8'h00}, /* 0xaaac */
            {8'h00}, /* 0xaaab */
            {8'h00}, /* 0xaaaa */
            {8'h00}, /* 0xaaa9 */
            {8'h00}, /* 0xaaa8 */
            {8'h00}, /* 0xaaa7 */
            {8'h00}, /* 0xaaa6 */
            {8'h00}, /* 0xaaa5 */
            {8'h00}, /* 0xaaa4 */
            {8'h00}, /* 0xaaa3 */
            {8'h00}, /* 0xaaa2 */
            {8'h00}, /* 0xaaa1 */
            {8'h00}, /* 0xaaa0 */
            {8'h00}, /* 0xaa9f */
            {8'h00}, /* 0xaa9e */
            {8'h00}, /* 0xaa9d */
            {8'h00}, /* 0xaa9c */
            {8'h00}, /* 0xaa9b */
            {8'h00}, /* 0xaa9a */
            {8'h00}, /* 0xaa99 */
            {8'h00}, /* 0xaa98 */
            {8'h00}, /* 0xaa97 */
            {8'h00}, /* 0xaa96 */
            {8'h00}, /* 0xaa95 */
            {8'h00}, /* 0xaa94 */
            {8'h00}, /* 0xaa93 */
            {8'h00}, /* 0xaa92 */
            {8'h00}, /* 0xaa91 */
            {8'h00}, /* 0xaa90 */
            {8'h00}, /* 0xaa8f */
            {8'h00}, /* 0xaa8e */
            {8'h00}, /* 0xaa8d */
            {8'h00}, /* 0xaa8c */
            {8'h00}, /* 0xaa8b */
            {8'h00}, /* 0xaa8a */
            {8'h00}, /* 0xaa89 */
            {8'h00}, /* 0xaa88 */
            {8'h00}, /* 0xaa87 */
            {8'h00}, /* 0xaa86 */
            {8'h00}, /* 0xaa85 */
            {8'h00}, /* 0xaa84 */
            {8'h00}, /* 0xaa83 */
            {8'h00}, /* 0xaa82 */
            {8'h00}, /* 0xaa81 */
            {8'h00}, /* 0xaa80 */
            {8'h00}, /* 0xaa7f */
            {8'h00}, /* 0xaa7e */
            {8'h00}, /* 0xaa7d */
            {8'h00}, /* 0xaa7c */
            {8'h00}, /* 0xaa7b */
            {8'h00}, /* 0xaa7a */
            {8'h00}, /* 0xaa79 */
            {8'h00}, /* 0xaa78 */
            {8'h00}, /* 0xaa77 */
            {8'h00}, /* 0xaa76 */
            {8'h00}, /* 0xaa75 */
            {8'h00}, /* 0xaa74 */
            {8'h00}, /* 0xaa73 */
            {8'h00}, /* 0xaa72 */
            {8'h00}, /* 0xaa71 */
            {8'h00}, /* 0xaa70 */
            {8'h00}, /* 0xaa6f */
            {8'h00}, /* 0xaa6e */
            {8'h00}, /* 0xaa6d */
            {8'h00}, /* 0xaa6c */
            {8'h00}, /* 0xaa6b */
            {8'h00}, /* 0xaa6a */
            {8'h00}, /* 0xaa69 */
            {8'h00}, /* 0xaa68 */
            {8'h00}, /* 0xaa67 */
            {8'h00}, /* 0xaa66 */
            {8'h00}, /* 0xaa65 */
            {8'h00}, /* 0xaa64 */
            {8'h00}, /* 0xaa63 */
            {8'h00}, /* 0xaa62 */
            {8'h00}, /* 0xaa61 */
            {8'h00}, /* 0xaa60 */
            {8'h00}, /* 0xaa5f */
            {8'h00}, /* 0xaa5e */
            {8'h00}, /* 0xaa5d */
            {8'h00}, /* 0xaa5c */
            {8'h00}, /* 0xaa5b */
            {8'h00}, /* 0xaa5a */
            {8'h00}, /* 0xaa59 */
            {8'h00}, /* 0xaa58 */
            {8'h00}, /* 0xaa57 */
            {8'h00}, /* 0xaa56 */
            {8'h00}, /* 0xaa55 */
            {8'h00}, /* 0xaa54 */
            {8'h00}, /* 0xaa53 */
            {8'h00}, /* 0xaa52 */
            {8'h00}, /* 0xaa51 */
            {8'h00}, /* 0xaa50 */
            {8'h00}, /* 0xaa4f */
            {8'h00}, /* 0xaa4e */
            {8'h00}, /* 0xaa4d */
            {8'h00}, /* 0xaa4c */
            {8'h00}, /* 0xaa4b */
            {8'h00}, /* 0xaa4a */
            {8'h00}, /* 0xaa49 */
            {8'h00}, /* 0xaa48 */
            {8'h00}, /* 0xaa47 */
            {8'h00}, /* 0xaa46 */
            {8'h00}, /* 0xaa45 */
            {8'h00}, /* 0xaa44 */
            {8'h00}, /* 0xaa43 */
            {8'h00}, /* 0xaa42 */
            {8'h00}, /* 0xaa41 */
            {8'h00}, /* 0xaa40 */
            {8'h00}, /* 0xaa3f */
            {8'h00}, /* 0xaa3e */
            {8'h00}, /* 0xaa3d */
            {8'h00}, /* 0xaa3c */
            {8'h00}, /* 0xaa3b */
            {8'h00}, /* 0xaa3a */
            {8'h00}, /* 0xaa39 */
            {8'h00}, /* 0xaa38 */
            {8'h00}, /* 0xaa37 */
            {8'h00}, /* 0xaa36 */
            {8'h00}, /* 0xaa35 */
            {8'h00}, /* 0xaa34 */
            {8'h00}, /* 0xaa33 */
            {8'h00}, /* 0xaa32 */
            {8'h00}, /* 0xaa31 */
            {8'h00}, /* 0xaa30 */
            {8'h00}, /* 0xaa2f */
            {8'h00}, /* 0xaa2e */
            {8'h00}, /* 0xaa2d */
            {8'h00}, /* 0xaa2c */
            {8'h00}, /* 0xaa2b */
            {8'h00}, /* 0xaa2a */
            {8'h00}, /* 0xaa29 */
            {8'h00}, /* 0xaa28 */
            {8'h00}, /* 0xaa27 */
            {8'h00}, /* 0xaa26 */
            {8'h00}, /* 0xaa25 */
            {8'h00}, /* 0xaa24 */
            {8'h00}, /* 0xaa23 */
            {8'h00}, /* 0xaa22 */
            {8'h00}, /* 0xaa21 */
            {8'h00}, /* 0xaa20 */
            {8'h00}, /* 0xaa1f */
            {8'h00}, /* 0xaa1e */
            {8'h00}, /* 0xaa1d */
            {8'h00}, /* 0xaa1c */
            {8'h00}, /* 0xaa1b */
            {8'h00}, /* 0xaa1a */
            {8'h00}, /* 0xaa19 */
            {8'h00}, /* 0xaa18 */
            {8'h00}, /* 0xaa17 */
            {8'h00}, /* 0xaa16 */
            {8'h00}, /* 0xaa15 */
            {8'h00}, /* 0xaa14 */
            {8'h00}, /* 0xaa13 */
            {8'h00}, /* 0xaa12 */
            {8'h00}, /* 0xaa11 */
            {8'h00}, /* 0xaa10 */
            {8'h00}, /* 0xaa0f */
            {8'h00}, /* 0xaa0e */
            {8'h00}, /* 0xaa0d */
            {8'h00}, /* 0xaa0c */
            {8'h00}, /* 0xaa0b */
            {8'h00}, /* 0xaa0a */
            {8'h00}, /* 0xaa09 */
            {8'h00}, /* 0xaa08 */
            {8'h00}, /* 0xaa07 */
            {8'h00}, /* 0xaa06 */
            {8'h00}, /* 0xaa05 */
            {8'h00}, /* 0xaa04 */
            {8'h00}, /* 0xaa03 */
            {8'h00}, /* 0xaa02 */
            {8'h00}, /* 0xaa01 */
            {8'h00}, /* 0xaa00 */
            {8'h00}, /* 0xa9ff */
            {8'h00}, /* 0xa9fe */
            {8'h00}, /* 0xa9fd */
            {8'h00}, /* 0xa9fc */
            {8'h00}, /* 0xa9fb */
            {8'h00}, /* 0xa9fa */
            {8'h00}, /* 0xa9f9 */
            {8'h00}, /* 0xa9f8 */
            {8'h00}, /* 0xa9f7 */
            {8'h00}, /* 0xa9f6 */
            {8'h00}, /* 0xa9f5 */
            {8'h00}, /* 0xa9f4 */
            {8'h00}, /* 0xa9f3 */
            {8'h00}, /* 0xa9f2 */
            {8'h00}, /* 0xa9f1 */
            {8'h00}, /* 0xa9f0 */
            {8'h00}, /* 0xa9ef */
            {8'h00}, /* 0xa9ee */
            {8'h00}, /* 0xa9ed */
            {8'h00}, /* 0xa9ec */
            {8'h00}, /* 0xa9eb */
            {8'h00}, /* 0xa9ea */
            {8'h00}, /* 0xa9e9 */
            {8'h00}, /* 0xa9e8 */
            {8'h00}, /* 0xa9e7 */
            {8'h00}, /* 0xa9e6 */
            {8'h00}, /* 0xa9e5 */
            {8'h00}, /* 0xa9e4 */
            {8'h00}, /* 0xa9e3 */
            {8'h00}, /* 0xa9e2 */
            {8'h00}, /* 0xa9e1 */
            {8'h00}, /* 0xa9e0 */
            {8'h00}, /* 0xa9df */
            {8'h00}, /* 0xa9de */
            {8'h00}, /* 0xa9dd */
            {8'h00}, /* 0xa9dc */
            {8'h00}, /* 0xa9db */
            {8'h00}, /* 0xa9da */
            {8'h00}, /* 0xa9d9 */
            {8'h00}, /* 0xa9d8 */
            {8'h00}, /* 0xa9d7 */
            {8'h00}, /* 0xa9d6 */
            {8'h00}, /* 0xa9d5 */
            {8'h00}, /* 0xa9d4 */
            {8'h00}, /* 0xa9d3 */
            {8'h00}, /* 0xa9d2 */
            {8'h00}, /* 0xa9d1 */
            {8'h00}, /* 0xa9d0 */
            {8'h00}, /* 0xa9cf */
            {8'h00}, /* 0xa9ce */
            {8'h00}, /* 0xa9cd */
            {8'h00}, /* 0xa9cc */
            {8'h00}, /* 0xa9cb */
            {8'h00}, /* 0xa9ca */
            {8'h00}, /* 0xa9c9 */
            {8'h00}, /* 0xa9c8 */
            {8'h00}, /* 0xa9c7 */
            {8'h00}, /* 0xa9c6 */
            {8'h00}, /* 0xa9c5 */
            {8'h00}, /* 0xa9c4 */
            {8'h00}, /* 0xa9c3 */
            {8'h00}, /* 0xa9c2 */
            {8'h00}, /* 0xa9c1 */
            {8'h00}, /* 0xa9c0 */
            {8'h00}, /* 0xa9bf */
            {8'h00}, /* 0xa9be */
            {8'h00}, /* 0xa9bd */
            {8'h00}, /* 0xa9bc */
            {8'h00}, /* 0xa9bb */
            {8'h00}, /* 0xa9ba */
            {8'h00}, /* 0xa9b9 */
            {8'h00}, /* 0xa9b8 */
            {8'h00}, /* 0xa9b7 */
            {8'h00}, /* 0xa9b6 */
            {8'h00}, /* 0xa9b5 */
            {8'h00}, /* 0xa9b4 */
            {8'h00}, /* 0xa9b3 */
            {8'h00}, /* 0xa9b2 */
            {8'h00}, /* 0xa9b1 */
            {8'h00}, /* 0xa9b0 */
            {8'h00}, /* 0xa9af */
            {8'h00}, /* 0xa9ae */
            {8'h00}, /* 0xa9ad */
            {8'h00}, /* 0xa9ac */
            {8'h00}, /* 0xa9ab */
            {8'h00}, /* 0xa9aa */
            {8'h00}, /* 0xa9a9 */
            {8'h00}, /* 0xa9a8 */
            {8'h00}, /* 0xa9a7 */
            {8'h00}, /* 0xa9a6 */
            {8'h00}, /* 0xa9a5 */
            {8'h00}, /* 0xa9a4 */
            {8'h00}, /* 0xa9a3 */
            {8'h00}, /* 0xa9a2 */
            {8'h00}, /* 0xa9a1 */
            {8'h00}, /* 0xa9a0 */
            {8'h00}, /* 0xa99f */
            {8'h00}, /* 0xa99e */
            {8'h00}, /* 0xa99d */
            {8'h00}, /* 0xa99c */
            {8'h00}, /* 0xa99b */
            {8'h00}, /* 0xa99a */
            {8'h00}, /* 0xa999 */
            {8'h00}, /* 0xa998 */
            {8'h00}, /* 0xa997 */
            {8'h00}, /* 0xa996 */
            {8'h00}, /* 0xa995 */
            {8'h00}, /* 0xa994 */
            {8'h00}, /* 0xa993 */
            {8'h00}, /* 0xa992 */
            {8'h00}, /* 0xa991 */
            {8'h00}, /* 0xa990 */
            {8'h00}, /* 0xa98f */
            {8'h00}, /* 0xa98e */
            {8'h00}, /* 0xa98d */
            {8'h00}, /* 0xa98c */
            {8'h00}, /* 0xa98b */
            {8'h00}, /* 0xa98a */
            {8'h00}, /* 0xa989 */
            {8'h00}, /* 0xa988 */
            {8'h00}, /* 0xa987 */
            {8'h00}, /* 0xa986 */
            {8'h00}, /* 0xa985 */
            {8'h00}, /* 0xa984 */
            {8'h00}, /* 0xa983 */
            {8'h00}, /* 0xa982 */
            {8'h00}, /* 0xa981 */
            {8'h00}, /* 0xa980 */
            {8'h00}, /* 0xa97f */
            {8'h00}, /* 0xa97e */
            {8'h00}, /* 0xa97d */
            {8'h00}, /* 0xa97c */
            {8'h00}, /* 0xa97b */
            {8'h00}, /* 0xa97a */
            {8'h00}, /* 0xa979 */
            {8'h00}, /* 0xa978 */
            {8'h00}, /* 0xa977 */
            {8'h00}, /* 0xa976 */
            {8'h00}, /* 0xa975 */
            {8'h00}, /* 0xa974 */
            {8'h00}, /* 0xa973 */
            {8'h00}, /* 0xa972 */
            {8'h00}, /* 0xa971 */
            {8'h00}, /* 0xa970 */
            {8'h00}, /* 0xa96f */
            {8'h00}, /* 0xa96e */
            {8'h00}, /* 0xa96d */
            {8'h00}, /* 0xa96c */
            {8'h00}, /* 0xa96b */
            {8'h00}, /* 0xa96a */
            {8'h00}, /* 0xa969 */
            {8'h00}, /* 0xa968 */
            {8'h00}, /* 0xa967 */
            {8'h00}, /* 0xa966 */
            {8'h00}, /* 0xa965 */
            {8'h00}, /* 0xa964 */
            {8'h00}, /* 0xa963 */
            {8'h00}, /* 0xa962 */
            {8'h00}, /* 0xa961 */
            {8'h00}, /* 0xa960 */
            {8'h00}, /* 0xa95f */
            {8'h00}, /* 0xa95e */
            {8'h00}, /* 0xa95d */
            {8'h00}, /* 0xa95c */
            {8'h00}, /* 0xa95b */
            {8'h00}, /* 0xa95a */
            {8'h00}, /* 0xa959 */
            {8'h00}, /* 0xa958 */
            {8'h00}, /* 0xa957 */
            {8'h00}, /* 0xa956 */
            {8'h00}, /* 0xa955 */
            {8'h00}, /* 0xa954 */
            {8'h00}, /* 0xa953 */
            {8'h00}, /* 0xa952 */
            {8'h00}, /* 0xa951 */
            {8'h00}, /* 0xa950 */
            {8'h00}, /* 0xa94f */
            {8'h00}, /* 0xa94e */
            {8'h00}, /* 0xa94d */
            {8'h00}, /* 0xa94c */
            {8'h00}, /* 0xa94b */
            {8'h00}, /* 0xa94a */
            {8'h00}, /* 0xa949 */
            {8'h00}, /* 0xa948 */
            {8'h00}, /* 0xa947 */
            {8'h00}, /* 0xa946 */
            {8'h00}, /* 0xa945 */
            {8'h00}, /* 0xa944 */
            {8'h00}, /* 0xa943 */
            {8'h00}, /* 0xa942 */
            {8'h00}, /* 0xa941 */
            {8'h00}, /* 0xa940 */
            {8'h00}, /* 0xa93f */
            {8'h00}, /* 0xa93e */
            {8'h00}, /* 0xa93d */
            {8'h00}, /* 0xa93c */
            {8'h00}, /* 0xa93b */
            {8'h00}, /* 0xa93a */
            {8'h00}, /* 0xa939 */
            {8'h00}, /* 0xa938 */
            {8'h00}, /* 0xa937 */
            {8'h00}, /* 0xa936 */
            {8'h00}, /* 0xa935 */
            {8'h00}, /* 0xa934 */
            {8'h00}, /* 0xa933 */
            {8'h00}, /* 0xa932 */
            {8'h00}, /* 0xa931 */
            {8'h00}, /* 0xa930 */
            {8'h00}, /* 0xa92f */
            {8'h00}, /* 0xa92e */
            {8'h00}, /* 0xa92d */
            {8'h00}, /* 0xa92c */
            {8'h00}, /* 0xa92b */
            {8'h00}, /* 0xa92a */
            {8'h00}, /* 0xa929 */
            {8'h00}, /* 0xa928 */
            {8'h00}, /* 0xa927 */
            {8'h00}, /* 0xa926 */
            {8'h00}, /* 0xa925 */
            {8'h00}, /* 0xa924 */
            {8'h00}, /* 0xa923 */
            {8'h00}, /* 0xa922 */
            {8'h00}, /* 0xa921 */
            {8'h00}, /* 0xa920 */
            {8'h00}, /* 0xa91f */
            {8'h00}, /* 0xa91e */
            {8'h00}, /* 0xa91d */
            {8'h00}, /* 0xa91c */
            {8'h00}, /* 0xa91b */
            {8'h00}, /* 0xa91a */
            {8'h00}, /* 0xa919 */
            {8'h00}, /* 0xa918 */
            {8'h00}, /* 0xa917 */
            {8'h00}, /* 0xa916 */
            {8'h00}, /* 0xa915 */
            {8'h00}, /* 0xa914 */
            {8'h00}, /* 0xa913 */
            {8'h00}, /* 0xa912 */
            {8'h00}, /* 0xa911 */
            {8'h00}, /* 0xa910 */
            {8'h00}, /* 0xa90f */
            {8'h00}, /* 0xa90e */
            {8'h00}, /* 0xa90d */
            {8'h00}, /* 0xa90c */
            {8'h00}, /* 0xa90b */
            {8'h00}, /* 0xa90a */
            {8'h00}, /* 0xa909 */
            {8'h00}, /* 0xa908 */
            {8'h00}, /* 0xa907 */
            {8'h00}, /* 0xa906 */
            {8'h00}, /* 0xa905 */
            {8'h00}, /* 0xa904 */
            {8'h00}, /* 0xa903 */
            {8'h00}, /* 0xa902 */
            {8'h00}, /* 0xa901 */
            {8'h00}, /* 0xa900 */
            {8'h00}, /* 0xa8ff */
            {8'h00}, /* 0xa8fe */
            {8'h00}, /* 0xa8fd */
            {8'h00}, /* 0xa8fc */
            {8'h00}, /* 0xa8fb */
            {8'h00}, /* 0xa8fa */
            {8'h00}, /* 0xa8f9 */
            {8'h00}, /* 0xa8f8 */
            {8'h00}, /* 0xa8f7 */
            {8'h00}, /* 0xa8f6 */
            {8'h00}, /* 0xa8f5 */
            {8'h00}, /* 0xa8f4 */
            {8'h00}, /* 0xa8f3 */
            {8'h00}, /* 0xa8f2 */
            {8'h00}, /* 0xa8f1 */
            {8'h00}, /* 0xa8f0 */
            {8'h00}, /* 0xa8ef */
            {8'h00}, /* 0xa8ee */
            {8'h00}, /* 0xa8ed */
            {8'h00}, /* 0xa8ec */
            {8'h00}, /* 0xa8eb */
            {8'h00}, /* 0xa8ea */
            {8'h00}, /* 0xa8e9 */
            {8'h00}, /* 0xa8e8 */
            {8'h00}, /* 0xa8e7 */
            {8'h00}, /* 0xa8e6 */
            {8'h00}, /* 0xa8e5 */
            {8'h00}, /* 0xa8e4 */
            {8'h00}, /* 0xa8e3 */
            {8'h00}, /* 0xa8e2 */
            {8'h00}, /* 0xa8e1 */
            {8'h00}, /* 0xa8e0 */
            {8'h00}, /* 0xa8df */
            {8'h00}, /* 0xa8de */
            {8'h00}, /* 0xa8dd */
            {8'h00}, /* 0xa8dc */
            {8'h00}, /* 0xa8db */
            {8'h00}, /* 0xa8da */
            {8'h00}, /* 0xa8d9 */
            {8'h00}, /* 0xa8d8 */
            {8'h00}, /* 0xa8d7 */
            {8'h00}, /* 0xa8d6 */
            {8'h00}, /* 0xa8d5 */
            {8'h00}, /* 0xa8d4 */
            {8'h00}, /* 0xa8d3 */
            {8'h00}, /* 0xa8d2 */
            {8'h00}, /* 0xa8d1 */
            {8'h00}, /* 0xa8d0 */
            {8'h00}, /* 0xa8cf */
            {8'h00}, /* 0xa8ce */
            {8'h00}, /* 0xa8cd */
            {8'h00}, /* 0xa8cc */
            {8'h00}, /* 0xa8cb */
            {8'h00}, /* 0xa8ca */
            {8'h00}, /* 0xa8c9 */
            {8'h00}, /* 0xa8c8 */
            {8'h00}, /* 0xa8c7 */
            {8'h00}, /* 0xa8c6 */
            {8'h00}, /* 0xa8c5 */
            {8'h00}, /* 0xa8c4 */
            {8'h00}, /* 0xa8c3 */
            {8'h00}, /* 0xa8c2 */
            {8'h00}, /* 0xa8c1 */
            {8'h00}, /* 0xa8c0 */
            {8'h00}, /* 0xa8bf */
            {8'h00}, /* 0xa8be */
            {8'h00}, /* 0xa8bd */
            {8'h00}, /* 0xa8bc */
            {8'h00}, /* 0xa8bb */
            {8'h00}, /* 0xa8ba */
            {8'h00}, /* 0xa8b9 */
            {8'h00}, /* 0xa8b8 */
            {8'h00}, /* 0xa8b7 */
            {8'h00}, /* 0xa8b6 */
            {8'h00}, /* 0xa8b5 */
            {8'h00}, /* 0xa8b4 */
            {8'h00}, /* 0xa8b3 */
            {8'h00}, /* 0xa8b2 */
            {8'h00}, /* 0xa8b1 */
            {8'h00}, /* 0xa8b0 */
            {8'h00}, /* 0xa8af */
            {8'h00}, /* 0xa8ae */
            {8'h00}, /* 0xa8ad */
            {8'h00}, /* 0xa8ac */
            {8'h00}, /* 0xa8ab */
            {8'h00}, /* 0xa8aa */
            {8'h00}, /* 0xa8a9 */
            {8'h00}, /* 0xa8a8 */
            {8'h00}, /* 0xa8a7 */
            {8'h00}, /* 0xa8a6 */
            {8'h00}, /* 0xa8a5 */
            {8'h00}, /* 0xa8a4 */
            {8'h00}, /* 0xa8a3 */
            {8'h00}, /* 0xa8a2 */
            {8'h00}, /* 0xa8a1 */
            {8'h00}, /* 0xa8a0 */
            {8'h00}, /* 0xa89f */
            {8'h00}, /* 0xa89e */
            {8'h00}, /* 0xa89d */
            {8'h00}, /* 0xa89c */
            {8'h00}, /* 0xa89b */
            {8'h00}, /* 0xa89a */
            {8'h00}, /* 0xa899 */
            {8'h00}, /* 0xa898 */
            {8'h00}, /* 0xa897 */
            {8'h00}, /* 0xa896 */
            {8'h00}, /* 0xa895 */
            {8'h00}, /* 0xa894 */
            {8'h00}, /* 0xa893 */
            {8'h00}, /* 0xa892 */
            {8'h00}, /* 0xa891 */
            {8'h00}, /* 0xa890 */
            {8'h00}, /* 0xa88f */
            {8'h00}, /* 0xa88e */
            {8'h00}, /* 0xa88d */
            {8'h00}, /* 0xa88c */
            {8'h00}, /* 0xa88b */
            {8'h00}, /* 0xa88a */
            {8'h00}, /* 0xa889 */
            {8'h00}, /* 0xa888 */
            {8'h00}, /* 0xa887 */
            {8'h00}, /* 0xa886 */
            {8'h00}, /* 0xa885 */
            {8'h00}, /* 0xa884 */
            {8'h00}, /* 0xa883 */
            {8'h00}, /* 0xa882 */
            {8'h00}, /* 0xa881 */
            {8'h00}, /* 0xa880 */
            {8'h00}, /* 0xa87f */
            {8'h00}, /* 0xa87e */
            {8'h00}, /* 0xa87d */
            {8'h00}, /* 0xa87c */
            {8'h00}, /* 0xa87b */
            {8'h00}, /* 0xa87a */
            {8'h00}, /* 0xa879 */
            {8'h00}, /* 0xa878 */
            {8'h00}, /* 0xa877 */
            {8'h00}, /* 0xa876 */
            {8'h00}, /* 0xa875 */
            {8'h00}, /* 0xa874 */
            {8'h00}, /* 0xa873 */
            {8'h00}, /* 0xa872 */
            {8'h00}, /* 0xa871 */
            {8'h00}, /* 0xa870 */
            {8'h00}, /* 0xa86f */
            {8'h00}, /* 0xa86e */
            {8'h00}, /* 0xa86d */
            {8'h00}, /* 0xa86c */
            {8'h00}, /* 0xa86b */
            {8'h00}, /* 0xa86a */
            {8'h00}, /* 0xa869 */
            {8'h00}, /* 0xa868 */
            {8'h00}, /* 0xa867 */
            {8'h00}, /* 0xa866 */
            {8'h00}, /* 0xa865 */
            {8'h00}, /* 0xa864 */
            {8'h00}, /* 0xa863 */
            {8'h00}, /* 0xa862 */
            {8'h00}, /* 0xa861 */
            {8'h00}, /* 0xa860 */
            {8'h00}, /* 0xa85f */
            {8'h00}, /* 0xa85e */
            {8'h00}, /* 0xa85d */
            {8'h00}, /* 0xa85c */
            {8'h00}, /* 0xa85b */
            {8'h00}, /* 0xa85a */
            {8'h00}, /* 0xa859 */
            {8'h00}, /* 0xa858 */
            {8'h00}, /* 0xa857 */
            {8'h00}, /* 0xa856 */
            {8'h00}, /* 0xa855 */
            {8'h00}, /* 0xa854 */
            {8'h00}, /* 0xa853 */
            {8'h00}, /* 0xa852 */
            {8'h00}, /* 0xa851 */
            {8'h00}, /* 0xa850 */
            {8'h00}, /* 0xa84f */
            {8'h00}, /* 0xa84e */
            {8'h00}, /* 0xa84d */
            {8'h00}, /* 0xa84c */
            {8'h00}, /* 0xa84b */
            {8'h00}, /* 0xa84a */
            {8'h00}, /* 0xa849 */
            {8'h00}, /* 0xa848 */
            {8'h00}, /* 0xa847 */
            {8'h00}, /* 0xa846 */
            {8'h00}, /* 0xa845 */
            {8'h00}, /* 0xa844 */
            {8'h00}, /* 0xa843 */
            {8'h00}, /* 0xa842 */
            {8'h00}, /* 0xa841 */
            {8'h00}, /* 0xa840 */
            {8'h00}, /* 0xa83f */
            {8'h00}, /* 0xa83e */
            {8'h00}, /* 0xa83d */
            {8'h00}, /* 0xa83c */
            {8'h00}, /* 0xa83b */
            {8'h00}, /* 0xa83a */
            {8'h00}, /* 0xa839 */
            {8'h00}, /* 0xa838 */
            {8'h00}, /* 0xa837 */
            {8'h00}, /* 0xa836 */
            {8'h00}, /* 0xa835 */
            {8'h00}, /* 0xa834 */
            {8'h00}, /* 0xa833 */
            {8'h00}, /* 0xa832 */
            {8'h00}, /* 0xa831 */
            {8'h00}, /* 0xa830 */
            {8'h00}, /* 0xa82f */
            {8'h00}, /* 0xa82e */
            {8'h00}, /* 0xa82d */
            {8'h00}, /* 0xa82c */
            {8'h00}, /* 0xa82b */
            {8'h00}, /* 0xa82a */
            {8'h00}, /* 0xa829 */
            {8'h00}, /* 0xa828 */
            {8'h00}, /* 0xa827 */
            {8'h00}, /* 0xa826 */
            {8'h00}, /* 0xa825 */
            {8'h00}, /* 0xa824 */
            {8'h00}, /* 0xa823 */
            {8'h00}, /* 0xa822 */
            {8'h00}, /* 0xa821 */
            {8'h00}, /* 0xa820 */
            {8'h00}, /* 0xa81f */
            {8'h00}, /* 0xa81e */
            {8'h00}, /* 0xa81d */
            {8'h00}, /* 0xa81c */
            {8'h00}, /* 0xa81b */
            {8'h00}, /* 0xa81a */
            {8'h00}, /* 0xa819 */
            {8'h00}, /* 0xa818 */
            {8'h00}, /* 0xa817 */
            {8'h00}, /* 0xa816 */
            {8'h00}, /* 0xa815 */
            {8'h00}, /* 0xa814 */
            {8'h00}, /* 0xa813 */
            {8'h00}, /* 0xa812 */
            {8'h00}, /* 0xa811 */
            {8'h00}, /* 0xa810 */
            {8'h00}, /* 0xa80f */
            {8'h00}, /* 0xa80e */
            {8'h00}, /* 0xa80d */
            {8'h00}, /* 0xa80c */
            {8'h00}, /* 0xa80b */
            {8'h00}, /* 0xa80a */
            {8'h00}, /* 0xa809 */
            {8'h00}, /* 0xa808 */
            {8'h00}, /* 0xa807 */
            {8'h00}, /* 0xa806 */
            {8'h00}, /* 0xa805 */
            {8'h00}, /* 0xa804 */
            {8'h00}, /* 0xa803 */
            {8'h00}, /* 0xa802 */
            {8'h00}, /* 0xa801 */
            {8'h00}, /* 0xa800 */
            {8'h00}, /* 0xa7ff */
            {8'h00}, /* 0xa7fe */
            {8'h00}, /* 0xa7fd */
            {8'h00}, /* 0xa7fc */
            {8'h00}, /* 0xa7fb */
            {8'h00}, /* 0xa7fa */
            {8'h00}, /* 0xa7f9 */
            {8'h00}, /* 0xa7f8 */
            {8'h00}, /* 0xa7f7 */
            {8'h00}, /* 0xa7f6 */
            {8'h00}, /* 0xa7f5 */
            {8'h00}, /* 0xa7f4 */
            {8'h00}, /* 0xa7f3 */
            {8'h00}, /* 0xa7f2 */
            {8'h00}, /* 0xa7f1 */
            {8'h00}, /* 0xa7f0 */
            {8'h00}, /* 0xa7ef */
            {8'h00}, /* 0xa7ee */
            {8'h00}, /* 0xa7ed */
            {8'h00}, /* 0xa7ec */
            {8'h00}, /* 0xa7eb */
            {8'h00}, /* 0xa7ea */
            {8'h00}, /* 0xa7e9 */
            {8'h00}, /* 0xa7e8 */
            {8'h00}, /* 0xa7e7 */
            {8'h00}, /* 0xa7e6 */
            {8'h00}, /* 0xa7e5 */
            {8'h00}, /* 0xa7e4 */
            {8'h00}, /* 0xa7e3 */
            {8'h00}, /* 0xa7e2 */
            {8'h00}, /* 0xa7e1 */
            {8'h00}, /* 0xa7e0 */
            {8'h00}, /* 0xa7df */
            {8'h00}, /* 0xa7de */
            {8'h00}, /* 0xa7dd */
            {8'h00}, /* 0xa7dc */
            {8'h00}, /* 0xa7db */
            {8'h00}, /* 0xa7da */
            {8'h00}, /* 0xa7d9 */
            {8'h00}, /* 0xa7d8 */
            {8'h00}, /* 0xa7d7 */
            {8'h00}, /* 0xa7d6 */
            {8'h00}, /* 0xa7d5 */
            {8'h00}, /* 0xa7d4 */
            {8'h00}, /* 0xa7d3 */
            {8'h00}, /* 0xa7d2 */
            {8'h00}, /* 0xa7d1 */
            {8'h00}, /* 0xa7d0 */
            {8'h00}, /* 0xa7cf */
            {8'h00}, /* 0xa7ce */
            {8'h00}, /* 0xa7cd */
            {8'h00}, /* 0xa7cc */
            {8'h00}, /* 0xa7cb */
            {8'h00}, /* 0xa7ca */
            {8'h00}, /* 0xa7c9 */
            {8'h00}, /* 0xa7c8 */
            {8'h00}, /* 0xa7c7 */
            {8'h00}, /* 0xa7c6 */
            {8'h00}, /* 0xa7c5 */
            {8'h00}, /* 0xa7c4 */
            {8'h00}, /* 0xa7c3 */
            {8'h00}, /* 0xa7c2 */
            {8'h00}, /* 0xa7c1 */
            {8'h00}, /* 0xa7c0 */
            {8'h00}, /* 0xa7bf */
            {8'h00}, /* 0xa7be */
            {8'h00}, /* 0xa7bd */
            {8'h00}, /* 0xa7bc */
            {8'h00}, /* 0xa7bb */
            {8'h00}, /* 0xa7ba */
            {8'h00}, /* 0xa7b9 */
            {8'h00}, /* 0xa7b8 */
            {8'h00}, /* 0xa7b7 */
            {8'h00}, /* 0xa7b6 */
            {8'h00}, /* 0xa7b5 */
            {8'h00}, /* 0xa7b4 */
            {8'h00}, /* 0xa7b3 */
            {8'h00}, /* 0xa7b2 */
            {8'h00}, /* 0xa7b1 */
            {8'h00}, /* 0xa7b0 */
            {8'h00}, /* 0xa7af */
            {8'h00}, /* 0xa7ae */
            {8'h00}, /* 0xa7ad */
            {8'h00}, /* 0xa7ac */
            {8'h00}, /* 0xa7ab */
            {8'h00}, /* 0xa7aa */
            {8'h00}, /* 0xa7a9 */
            {8'h00}, /* 0xa7a8 */
            {8'h00}, /* 0xa7a7 */
            {8'h00}, /* 0xa7a6 */
            {8'h00}, /* 0xa7a5 */
            {8'h00}, /* 0xa7a4 */
            {8'h00}, /* 0xa7a3 */
            {8'h00}, /* 0xa7a2 */
            {8'h00}, /* 0xa7a1 */
            {8'h00}, /* 0xa7a0 */
            {8'h00}, /* 0xa79f */
            {8'h00}, /* 0xa79e */
            {8'h00}, /* 0xa79d */
            {8'h00}, /* 0xa79c */
            {8'h00}, /* 0xa79b */
            {8'h00}, /* 0xa79a */
            {8'h00}, /* 0xa799 */
            {8'h00}, /* 0xa798 */
            {8'h00}, /* 0xa797 */
            {8'h00}, /* 0xa796 */
            {8'h00}, /* 0xa795 */
            {8'h00}, /* 0xa794 */
            {8'h00}, /* 0xa793 */
            {8'h00}, /* 0xa792 */
            {8'h00}, /* 0xa791 */
            {8'h00}, /* 0xa790 */
            {8'h00}, /* 0xa78f */
            {8'h00}, /* 0xa78e */
            {8'h00}, /* 0xa78d */
            {8'h00}, /* 0xa78c */
            {8'h00}, /* 0xa78b */
            {8'h00}, /* 0xa78a */
            {8'h00}, /* 0xa789 */
            {8'h00}, /* 0xa788 */
            {8'h00}, /* 0xa787 */
            {8'h00}, /* 0xa786 */
            {8'h00}, /* 0xa785 */
            {8'h00}, /* 0xa784 */
            {8'h00}, /* 0xa783 */
            {8'h00}, /* 0xa782 */
            {8'h00}, /* 0xa781 */
            {8'h00}, /* 0xa780 */
            {8'h00}, /* 0xa77f */
            {8'h00}, /* 0xa77e */
            {8'h00}, /* 0xa77d */
            {8'h00}, /* 0xa77c */
            {8'h00}, /* 0xa77b */
            {8'h00}, /* 0xa77a */
            {8'h00}, /* 0xa779 */
            {8'h00}, /* 0xa778 */
            {8'h00}, /* 0xa777 */
            {8'h00}, /* 0xa776 */
            {8'h00}, /* 0xa775 */
            {8'h00}, /* 0xa774 */
            {8'h00}, /* 0xa773 */
            {8'h00}, /* 0xa772 */
            {8'h00}, /* 0xa771 */
            {8'h00}, /* 0xa770 */
            {8'h00}, /* 0xa76f */
            {8'h00}, /* 0xa76e */
            {8'h00}, /* 0xa76d */
            {8'h00}, /* 0xa76c */
            {8'h00}, /* 0xa76b */
            {8'h00}, /* 0xa76a */
            {8'h00}, /* 0xa769 */
            {8'h00}, /* 0xa768 */
            {8'h00}, /* 0xa767 */
            {8'h00}, /* 0xa766 */
            {8'h00}, /* 0xa765 */
            {8'h00}, /* 0xa764 */
            {8'h00}, /* 0xa763 */
            {8'h00}, /* 0xa762 */
            {8'h00}, /* 0xa761 */
            {8'h00}, /* 0xa760 */
            {8'h00}, /* 0xa75f */
            {8'h00}, /* 0xa75e */
            {8'h00}, /* 0xa75d */
            {8'h00}, /* 0xa75c */
            {8'h00}, /* 0xa75b */
            {8'h00}, /* 0xa75a */
            {8'h00}, /* 0xa759 */
            {8'h00}, /* 0xa758 */
            {8'h00}, /* 0xa757 */
            {8'h00}, /* 0xa756 */
            {8'h00}, /* 0xa755 */
            {8'h00}, /* 0xa754 */
            {8'h00}, /* 0xa753 */
            {8'h00}, /* 0xa752 */
            {8'h00}, /* 0xa751 */
            {8'h00}, /* 0xa750 */
            {8'h00}, /* 0xa74f */
            {8'h00}, /* 0xa74e */
            {8'h00}, /* 0xa74d */
            {8'h00}, /* 0xa74c */
            {8'h00}, /* 0xa74b */
            {8'h00}, /* 0xa74a */
            {8'h00}, /* 0xa749 */
            {8'h00}, /* 0xa748 */
            {8'h00}, /* 0xa747 */
            {8'h00}, /* 0xa746 */
            {8'h00}, /* 0xa745 */
            {8'h00}, /* 0xa744 */
            {8'h00}, /* 0xa743 */
            {8'h00}, /* 0xa742 */
            {8'h00}, /* 0xa741 */
            {8'h00}, /* 0xa740 */
            {8'h00}, /* 0xa73f */
            {8'h00}, /* 0xa73e */
            {8'h00}, /* 0xa73d */
            {8'h00}, /* 0xa73c */
            {8'h00}, /* 0xa73b */
            {8'h00}, /* 0xa73a */
            {8'h00}, /* 0xa739 */
            {8'h00}, /* 0xa738 */
            {8'h00}, /* 0xa737 */
            {8'h00}, /* 0xa736 */
            {8'h00}, /* 0xa735 */
            {8'h00}, /* 0xa734 */
            {8'h00}, /* 0xa733 */
            {8'h00}, /* 0xa732 */
            {8'h00}, /* 0xa731 */
            {8'h00}, /* 0xa730 */
            {8'h00}, /* 0xa72f */
            {8'h00}, /* 0xa72e */
            {8'h00}, /* 0xa72d */
            {8'h00}, /* 0xa72c */
            {8'h00}, /* 0xa72b */
            {8'h00}, /* 0xa72a */
            {8'h00}, /* 0xa729 */
            {8'h00}, /* 0xa728 */
            {8'h00}, /* 0xa727 */
            {8'h00}, /* 0xa726 */
            {8'h00}, /* 0xa725 */
            {8'h00}, /* 0xa724 */
            {8'h00}, /* 0xa723 */
            {8'h00}, /* 0xa722 */
            {8'h00}, /* 0xa721 */
            {8'h00}, /* 0xa720 */
            {8'h00}, /* 0xa71f */
            {8'h00}, /* 0xa71e */
            {8'h00}, /* 0xa71d */
            {8'h00}, /* 0xa71c */
            {8'h00}, /* 0xa71b */
            {8'h00}, /* 0xa71a */
            {8'h00}, /* 0xa719 */
            {8'h00}, /* 0xa718 */
            {8'h00}, /* 0xa717 */
            {8'h00}, /* 0xa716 */
            {8'h00}, /* 0xa715 */
            {8'h00}, /* 0xa714 */
            {8'h00}, /* 0xa713 */
            {8'h00}, /* 0xa712 */
            {8'h00}, /* 0xa711 */
            {8'h00}, /* 0xa710 */
            {8'h00}, /* 0xa70f */
            {8'h00}, /* 0xa70e */
            {8'h00}, /* 0xa70d */
            {8'h00}, /* 0xa70c */
            {8'h00}, /* 0xa70b */
            {8'h00}, /* 0xa70a */
            {8'h00}, /* 0xa709 */
            {8'h00}, /* 0xa708 */
            {8'h00}, /* 0xa707 */
            {8'h00}, /* 0xa706 */
            {8'h00}, /* 0xa705 */
            {8'h00}, /* 0xa704 */
            {8'h00}, /* 0xa703 */
            {8'h00}, /* 0xa702 */
            {8'h00}, /* 0xa701 */
            {8'h00}, /* 0xa700 */
            {8'h00}, /* 0xa6ff */
            {8'h00}, /* 0xa6fe */
            {8'h00}, /* 0xa6fd */
            {8'h00}, /* 0xa6fc */
            {8'h00}, /* 0xa6fb */
            {8'h00}, /* 0xa6fa */
            {8'h00}, /* 0xa6f9 */
            {8'h00}, /* 0xa6f8 */
            {8'h00}, /* 0xa6f7 */
            {8'h00}, /* 0xa6f6 */
            {8'h00}, /* 0xa6f5 */
            {8'h00}, /* 0xa6f4 */
            {8'h00}, /* 0xa6f3 */
            {8'h00}, /* 0xa6f2 */
            {8'h00}, /* 0xa6f1 */
            {8'h00}, /* 0xa6f0 */
            {8'h00}, /* 0xa6ef */
            {8'h00}, /* 0xa6ee */
            {8'h00}, /* 0xa6ed */
            {8'h00}, /* 0xa6ec */
            {8'h00}, /* 0xa6eb */
            {8'h00}, /* 0xa6ea */
            {8'h00}, /* 0xa6e9 */
            {8'h00}, /* 0xa6e8 */
            {8'h00}, /* 0xa6e7 */
            {8'h00}, /* 0xa6e6 */
            {8'h00}, /* 0xa6e5 */
            {8'h00}, /* 0xa6e4 */
            {8'h00}, /* 0xa6e3 */
            {8'h00}, /* 0xa6e2 */
            {8'h00}, /* 0xa6e1 */
            {8'h00}, /* 0xa6e0 */
            {8'h00}, /* 0xa6df */
            {8'h00}, /* 0xa6de */
            {8'h00}, /* 0xa6dd */
            {8'h00}, /* 0xa6dc */
            {8'h00}, /* 0xa6db */
            {8'h00}, /* 0xa6da */
            {8'h00}, /* 0xa6d9 */
            {8'h00}, /* 0xa6d8 */
            {8'h00}, /* 0xa6d7 */
            {8'h00}, /* 0xa6d6 */
            {8'h00}, /* 0xa6d5 */
            {8'h00}, /* 0xa6d4 */
            {8'h00}, /* 0xa6d3 */
            {8'h00}, /* 0xa6d2 */
            {8'h00}, /* 0xa6d1 */
            {8'h00}, /* 0xa6d0 */
            {8'h00}, /* 0xa6cf */
            {8'h00}, /* 0xa6ce */
            {8'h00}, /* 0xa6cd */
            {8'h00}, /* 0xa6cc */
            {8'h00}, /* 0xa6cb */
            {8'h00}, /* 0xa6ca */
            {8'h00}, /* 0xa6c9 */
            {8'h00}, /* 0xa6c8 */
            {8'h00}, /* 0xa6c7 */
            {8'h00}, /* 0xa6c6 */
            {8'h00}, /* 0xa6c5 */
            {8'h00}, /* 0xa6c4 */
            {8'h00}, /* 0xa6c3 */
            {8'h00}, /* 0xa6c2 */
            {8'h00}, /* 0xa6c1 */
            {8'h00}, /* 0xa6c0 */
            {8'h00}, /* 0xa6bf */
            {8'h00}, /* 0xa6be */
            {8'h00}, /* 0xa6bd */
            {8'h00}, /* 0xa6bc */
            {8'h00}, /* 0xa6bb */
            {8'h00}, /* 0xa6ba */
            {8'h00}, /* 0xa6b9 */
            {8'h00}, /* 0xa6b8 */
            {8'h00}, /* 0xa6b7 */
            {8'h00}, /* 0xa6b6 */
            {8'h00}, /* 0xa6b5 */
            {8'h00}, /* 0xa6b4 */
            {8'h00}, /* 0xa6b3 */
            {8'h00}, /* 0xa6b2 */
            {8'h00}, /* 0xa6b1 */
            {8'h00}, /* 0xa6b0 */
            {8'h00}, /* 0xa6af */
            {8'h00}, /* 0xa6ae */
            {8'h00}, /* 0xa6ad */
            {8'h00}, /* 0xa6ac */
            {8'h00}, /* 0xa6ab */
            {8'h00}, /* 0xa6aa */
            {8'h00}, /* 0xa6a9 */
            {8'h00}, /* 0xa6a8 */
            {8'h00}, /* 0xa6a7 */
            {8'h00}, /* 0xa6a6 */
            {8'h00}, /* 0xa6a5 */
            {8'h00}, /* 0xa6a4 */
            {8'h00}, /* 0xa6a3 */
            {8'h00}, /* 0xa6a2 */
            {8'h00}, /* 0xa6a1 */
            {8'h00}, /* 0xa6a0 */
            {8'h00}, /* 0xa69f */
            {8'h00}, /* 0xa69e */
            {8'h00}, /* 0xa69d */
            {8'h00}, /* 0xa69c */
            {8'h00}, /* 0xa69b */
            {8'h00}, /* 0xa69a */
            {8'h00}, /* 0xa699 */
            {8'h00}, /* 0xa698 */
            {8'h00}, /* 0xa697 */
            {8'h00}, /* 0xa696 */
            {8'h00}, /* 0xa695 */
            {8'h00}, /* 0xa694 */
            {8'h00}, /* 0xa693 */
            {8'h00}, /* 0xa692 */
            {8'h00}, /* 0xa691 */
            {8'h00}, /* 0xa690 */
            {8'h00}, /* 0xa68f */
            {8'h00}, /* 0xa68e */
            {8'h00}, /* 0xa68d */
            {8'h00}, /* 0xa68c */
            {8'h00}, /* 0xa68b */
            {8'h00}, /* 0xa68a */
            {8'h00}, /* 0xa689 */
            {8'h00}, /* 0xa688 */
            {8'h00}, /* 0xa687 */
            {8'h00}, /* 0xa686 */
            {8'h00}, /* 0xa685 */
            {8'h00}, /* 0xa684 */
            {8'h00}, /* 0xa683 */
            {8'h00}, /* 0xa682 */
            {8'h00}, /* 0xa681 */
            {8'h00}, /* 0xa680 */
            {8'h00}, /* 0xa67f */
            {8'h00}, /* 0xa67e */
            {8'h00}, /* 0xa67d */
            {8'h00}, /* 0xa67c */
            {8'h00}, /* 0xa67b */
            {8'h00}, /* 0xa67a */
            {8'h00}, /* 0xa679 */
            {8'h00}, /* 0xa678 */
            {8'h00}, /* 0xa677 */
            {8'h00}, /* 0xa676 */
            {8'h00}, /* 0xa675 */
            {8'h00}, /* 0xa674 */
            {8'h00}, /* 0xa673 */
            {8'h00}, /* 0xa672 */
            {8'h00}, /* 0xa671 */
            {8'h00}, /* 0xa670 */
            {8'h00}, /* 0xa66f */
            {8'h00}, /* 0xa66e */
            {8'h00}, /* 0xa66d */
            {8'h00}, /* 0xa66c */
            {8'h00}, /* 0xa66b */
            {8'h00}, /* 0xa66a */
            {8'h00}, /* 0xa669 */
            {8'h00}, /* 0xa668 */
            {8'h00}, /* 0xa667 */
            {8'h00}, /* 0xa666 */
            {8'h00}, /* 0xa665 */
            {8'h00}, /* 0xa664 */
            {8'h00}, /* 0xa663 */
            {8'h00}, /* 0xa662 */
            {8'h00}, /* 0xa661 */
            {8'h00}, /* 0xa660 */
            {8'h00}, /* 0xa65f */
            {8'h00}, /* 0xa65e */
            {8'h00}, /* 0xa65d */
            {8'h00}, /* 0xa65c */
            {8'h00}, /* 0xa65b */
            {8'h00}, /* 0xa65a */
            {8'h00}, /* 0xa659 */
            {8'h00}, /* 0xa658 */
            {8'h00}, /* 0xa657 */
            {8'h00}, /* 0xa656 */
            {8'h00}, /* 0xa655 */
            {8'h00}, /* 0xa654 */
            {8'h00}, /* 0xa653 */
            {8'h00}, /* 0xa652 */
            {8'h00}, /* 0xa651 */
            {8'h00}, /* 0xa650 */
            {8'h00}, /* 0xa64f */
            {8'h00}, /* 0xa64e */
            {8'h00}, /* 0xa64d */
            {8'h00}, /* 0xa64c */
            {8'h00}, /* 0xa64b */
            {8'h00}, /* 0xa64a */
            {8'h00}, /* 0xa649 */
            {8'h00}, /* 0xa648 */
            {8'h00}, /* 0xa647 */
            {8'h00}, /* 0xa646 */
            {8'h00}, /* 0xa645 */
            {8'h00}, /* 0xa644 */
            {8'h00}, /* 0xa643 */
            {8'h00}, /* 0xa642 */
            {8'h00}, /* 0xa641 */
            {8'h00}, /* 0xa640 */
            {8'h00}, /* 0xa63f */
            {8'h00}, /* 0xa63e */
            {8'h00}, /* 0xa63d */
            {8'h00}, /* 0xa63c */
            {8'h00}, /* 0xa63b */
            {8'h00}, /* 0xa63a */
            {8'h00}, /* 0xa639 */
            {8'h00}, /* 0xa638 */
            {8'h00}, /* 0xa637 */
            {8'h00}, /* 0xa636 */
            {8'h00}, /* 0xa635 */
            {8'h00}, /* 0xa634 */
            {8'h00}, /* 0xa633 */
            {8'h00}, /* 0xa632 */
            {8'h00}, /* 0xa631 */
            {8'h00}, /* 0xa630 */
            {8'h00}, /* 0xa62f */
            {8'h00}, /* 0xa62e */
            {8'h00}, /* 0xa62d */
            {8'h00}, /* 0xa62c */
            {8'h00}, /* 0xa62b */
            {8'h00}, /* 0xa62a */
            {8'h00}, /* 0xa629 */
            {8'h00}, /* 0xa628 */
            {8'h00}, /* 0xa627 */
            {8'h00}, /* 0xa626 */
            {8'h00}, /* 0xa625 */
            {8'h00}, /* 0xa624 */
            {8'h00}, /* 0xa623 */
            {8'h00}, /* 0xa622 */
            {8'h00}, /* 0xa621 */
            {8'h00}, /* 0xa620 */
            {8'h00}, /* 0xa61f */
            {8'h00}, /* 0xa61e */
            {8'h00}, /* 0xa61d */
            {8'h00}, /* 0xa61c */
            {8'h00}, /* 0xa61b */
            {8'h00}, /* 0xa61a */
            {8'h00}, /* 0xa619 */
            {8'h00}, /* 0xa618 */
            {8'h00}, /* 0xa617 */
            {8'h00}, /* 0xa616 */
            {8'h00}, /* 0xa615 */
            {8'h00}, /* 0xa614 */
            {8'h00}, /* 0xa613 */
            {8'h00}, /* 0xa612 */
            {8'h00}, /* 0xa611 */
            {8'h00}, /* 0xa610 */
            {8'h00}, /* 0xa60f */
            {8'h00}, /* 0xa60e */
            {8'h00}, /* 0xa60d */
            {8'h00}, /* 0xa60c */
            {8'h00}, /* 0xa60b */
            {8'h00}, /* 0xa60a */
            {8'h00}, /* 0xa609 */
            {8'h00}, /* 0xa608 */
            {8'h00}, /* 0xa607 */
            {8'h00}, /* 0xa606 */
            {8'h00}, /* 0xa605 */
            {8'h00}, /* 0xa604 */
            {8'h00}, /* 0xa603 */
            {8'h00}, /* 0xa602 */
            {8'h00}, /* 0xa601 */
            {8'h00}, /* 0xa600 */
            {8'h00}, /* 0xa5ff */
            {8'h00}, /* 0xa5fe */
            {8'h00}, /* 0xa5fd */
            {8'h00}, /* 0xa5fc */
            {8'h00}, /* 0xa5fb */
            {8'h00}, /* 0xa5fa */
            {8'h00}, /* 0xa5f9 */
            {8'h00}, /* 0xa5f8 */
            {8'h00}, /* 0xa5f7 */
            {8'h00}, /* 0xa5f6 */
            {8'h00}, /* 0xa5f5 */
            {8'h00}, /* 0xa5f4 */
            {8'h00}, /* 0xa5f3 */
            {8'h00}, /* 0xa5f2 */
            {8'h00}, /* 0xa5f1 */
            {8'h00}, /* 0xa5f0 */
            {8'h00}, /* 0xa5ef */
            {8'h00}, /* 0xa5ee */
            {8'h00}, /* 0xa5ed */
            {8'h00}, /* 0xa5ec */
            {8'h00}, /* 0xa5eb */
            {8'h00}, /* 0xa5ea */
            {8'h00}, /* 0xa5e9 */
            {8'h00}, /* 0xa5e8 */
            {8'h00}, /* 0xa5e7 */
            {8'h00}, /* 0xa5e6 */
            {8'h00}, /* 0xa5e5 */
            {8'h00}, /* 0xa5e4 */
            {8'h00}, /* 0xa5e3 */
            {8'h00}, /* 0xa5e2 */
            {8'h00}, /* 0xa5e1 */
            {8'h00}, /* 0xa5e0 */
            {8'h00}, /* 0xa5df */
            {8'h00}, /* 0xa5de */
            {8'h00}, /* 0xa5dd */
            {8'h00}, /* 0xa5dc */
            {8'h00}, /* 0xa5db */
            {8'h00}, /* 0xa5da */
            {8'h00}, /* 0xa5d9 */
            {8'h00}, /* 0xa5d8 */
            {8'h00}, /* 0xa5d7 */
            {8'h00}, /* 0xa5d6 */
            {8'h00}, /* 0xa5d5 */
            {8'h00}, /* 0xa5d4 */
            {8'h00}, /* 0xa5d3 */
            {8'h00}, /* 0xa5d2 */
            {8'h00}, /* 0xa5d1 */
            {8'h00}, /* 0xa5d0 */
            {8'h00}, /* 0xa5cf */
            {8'h00}, /* 0xa5ce */
            {8'h00}, /* 0xa5cd */
            {8'h00}, /* 0xa5cc */
            {8'h00}, /* 0xa5cb */
            {8'h00}, /* 0xa5ca */
            {8'h00}, /* 0xa5c9 */
            {8'h00}, /* 0xa5c8 */
            {8'h00}, /* 0xa5c7 */
            {8'h00}, /* 0xa5c6 */
            {8'h00}, /* 0xa5c5 */
            {8'h00}, /* 0xa5c4 */
            {8'h00}, /* 0xa5c3 */
            {8'h00}, /* 0xa5c2 */
            {8'h00}, /* 0xa5c1 */
            {8'h00}, /* 0xa5c0 */
            {8'h00}, /* 0xa5bf */
            {8'h00}, /* 0xa5be */
            {8'h00}, /* 0xa5bd */
            {8'h00}, /* 0xa5bc */
            {8'h00}, /* 0xa5bb */
            {8'h00}, /* 0xa5ba */
            {8'h00}, /* 0xa5b9 */
            {8'h00}, /* 0xa5b8 */
            {8'h00}, /* 0xa5b7 */
            {8'h00}, /* 0xa5b6 */
            {8'h00}, /* 0xa5b5 */
            {8'h00}, /* 0xa5b4 */
            {8'h00}, /* 0xa5b3 */
            {8'h00}, /* 0xa5b2 */
            {8'h00}, /* 0xa5b1 */
            {8'h00}, /* 0xa5b0 */
            {8'h00}, /* 0xa5af */
            {8'h00}, /* 0xa5ae */
            {8'h00}, /* 0xa5ad */
            {8'h00}, /* 0xa5ac */
            {8'h00}, /* 0xa5ab */
            {8'h00}, /* 0xa5aa */
            {8'h00}, /* 0xa5a9 */
            {8'h00}, /* 0xa5a8 */
            {8'h00}, /* 0xa5a7 */
            {8'h00}, /* 0xa5a6 */
            {8'h00}, /* 0xa5a5 */
            {8'h00}, /* 0xa5a4 */
            {8'h00}, /* 0xa5a3 */
            {8'h00}, /* 0xa5a2 */
            {8'h00}, /* 0xa5a1 */
            {8'h00}, /* 0xa5a0 */
            {8'h00}, /* 0xa59f */
            {8'h00}, /* 0xa59e */
            {8'h00}, /* 0xa59d */
            {8'h00}, /* 0xa59c */
            {8'h00}, /* 0xa59b */
            {8'h00}, /* 0xa59a */
            {8'h00}, /* 0xa599 */
            {8'h00}, /* 0xa598 */
            {8'h00}, /* 0xa597 */
            {8'h00}, /* 0xa596 */
            {8'h00}, /* 0xa595 */
            {8'h00}, /* 0xa594 */
            {8'h00}, /* 0xa593 */
            {8'h00}, /* 0xa592 */
            {8'h00}, /* 0xa591 */
            {8'h00}, /* 0xa590 */
            {8'h00}, /* 0xa58f */
            {8'h00}, /* 0xa58e */
            {8'h00}, /* 0xa58d */
            {8'h00}, /* 0xa58c */
            {8'h00}, /* 0xa58b */
            {8'h00}, /* 0xa58a */
            {8'h00}, /* 0xa589 */
            {8'h00}, /* 0xa588 */
            {8'h00}, /* 0xa587 */
            {8'h00}, /* 0xa586 */
            {8'h00}, /* 0xa585 */
            {8'h00}, /* 0xa584 */
            {8'h00}, /* 0xa583 */
            {8'h00}, /* 0xa582 */
            {8'h00}, /* 0xa581 */
            {8'h00}, /* 0xa580 */
            {8'h00}, /* 0xa57f */
            {8'h00}, /* 0xa57e */
            {8'h00}, /* 0xa57d */
            {8'h00}, /* 0xa57c */
            {8'h00}, /* 0xa57b */
            {8'h00}, /* 0xa57a */
            {8'h00}, /* 0xa579 */
            {8'h00}, /* 0xa578 */
            {8'h00}, /* 0xa577 */
            {8'h00}, /* 0xa576 */
            {8'h00}, /* 0xa575 */
            {8'h00}, /* 0xa574 */
            {8'h00}, /* 0xa573 */
            {8'h00}, /* 0xa572 */
            {8'h00}, /* 0xa571 */
            {8'h00}, /* 0xa570 */
            {8'h00}, /* 0xa56f */
            {8'h00}, /* 0xa56e */
            {8'h00}, /* 0xa56d */
            {8'h00}, /* 0xa56c */
            {8'h00}, /* 0xa56b */
            {8'h00}, /* 0xa56a */
            {8'h00}, /* 0xa569 */
            {8'h00}, /* 0xa568 */
            {8'h00}, /* 0xa567 */
            {8'h00}, /* 0xa566 */
            {8'h00}, /* 0xa565 */
            {8'h00}, /* 0xa564 */
            {8'h00}, /* 0xa563 */
            {8'h00}, /* 0xa562 */
            {8'h00}, /* 0xa561 */
            {8'h00}, /* 0xa560 */
            {8'h00}, /* 0xa55f */
            {8'h00}, /* 0xa55e */
            {8'h00}, /* 0xa55d */
            {8'h00}, /* 0xa55c */
            {8'h00}, /* 0xa55b */
            {8'h00}, /* 0xa55a */
            {8'h00}, /* 0xa559 */
            {8'h00}, /* 0xa558 */
            {8'h00}, /* 0xa557 */
            {8'h00}, /* 0xa556 */
            {8'h00}, /* 0xa555 */
            {8'h00}, /* 0xa554 */
            {8'h00}, /* 0xa553 */
            {8'h00}, /* 0xa552 */
            {8'h00}, /* 0xa551 */
            {8'h00}, /* 0xa550 */
            {8'h00}, /* 0xa54f */
            {8'h00}, /* 0xa54e */
            {8'h00}, /* 0xa54d */
            {8'h00}, /* 0xa54c */
            {8'h00}, /* 0xa54b */
            {8'h00}, /* 0xa54a */
            {8'h00}, /* 0xa549 */
            {8'h00}, /* 0xa548 */
            {8'h00}, /* 0xa547 */
            {8'h00}, /* 0xa546 */
            {8'h00}, /* 0xa545 */
            {8'h00}, /* 0xa544 */
            {8'h00}, /* 0xa543 */
            {8'h00}, /* 0xa542 */
            {8'h00}, /* 0xa541 */
            {8'h00}, /* 0xa540 */
            {8'h00}, /* 0xa53f */
            {8'h00}, /* 0xa53e */
            {8'h00}, /* 0xa53d */
            {8'h00}, /* 0xa53c */
            {8'h00}, /* 0xa53b */
            {8'h00}, /* 0xa53a */
            {8'h00}, /* 0xa539 */
            {8'h00}, /* 0xa538 */
            {8'h00}, /* 0xa537 */
            {8'h00}, /* 0xa536 */
            {8'h00}, /* 0xa535 */
            {8'h00}, /* 0xa534 */
            {8'h00}, /* 0xa533 */
            {8'h00}, /* 0xa532 */
            {8'h00}, /* 0xa531 */
            {8'h00}, /* 0xa530 */
            {8'h00}, /* 0xa52f */
            {8'h00}, /* 0xa52e */
            {8'h00}, /* 0xa52d */
            {8'h00}, /* 0xa52c */
            {8'h00}, /* 0xa52b */
            {8'h00}, /* 0xa52a */
            {8'h00}, /* 0xa529 */
            {8'h00}, /* 0xa528 */
            {8'h00}, /* 0xa527 */
            {8'h00}, /* 0xa526 */
            {8'h00}, /* 0xa525 */
            {8'h00}, /* 0xa524 */
            {8'h00}, /* 0xa523 */
            {8'h00}, /* 0xa522 */
            {8'h00}, /* 0xa521 */
            {8'h00}, /* 0xa520 */
            {8'h00}, /* 0xa51f */
            {8'h00}, /* 0xa51e */
            {8'h00}, /* 0xa51d */
            {8'h00}, /* 0xa51c */
            {8'h00}, /* 0xa51b */
            {8'h00}, /* 0xa51a */
            {8'h00}, /* 0xa519 */
            {8'h00}, /* 0xa518 */
            {8'h00}, /* 0xa517 */
            {8'h00}, /* 0xa516 */
            {8'h00}, /* 0xa515 */
            {8'h00}, /* 0xa514 */
            {8'h00}, /* 0xa513 */
            {8'h00}, /* 0xa512 */
            {8'h00}, /* 0xa511 */
            {8'h00}, /* 0xa510 */
            {8'h00}, /* 0xa50f */
            {8'h00}, /* 0xa50e */
            {8'h00}, /* 0xa50d */
            {8'h00}, /* 0xa50c */
            {8'h00}, /* 0xa50b */
            {8'h00}, /* 0xa50a */
            {8'h00}, /* 0xa509 */
            {8'h00}, /* 0xa508 */
            {8'h00}, /* 0xa507 */
            {8'h00}, /* 0xa506 */
            {8'h00}, /* 0xa505 */
            {8'h00}, /* 0xa504 */
            {8'h00}, /* 0xa503 */
            {8'h00}, /* 0xa502 */
            {8'h00}, /* 0xa501 */
            {8'h00}, /* 0xa500 */
            {8'h00}, /* 0xa4ff */
            {8'h00}, /* 0xa4fe */
            {8'h00}, /* 0xa4fd */
            {8'h00}, /* 0xa4fc */
            {8'h00}, /* 0xa4fb */
            {8'h00}, /* 0xa4fa */
            {8'h00}, /* 0xa4f9 */
            {8'h00}, /* 0xa4f8 */
            {8'h00}, /* 0xa4f7 */
            {8'h00}, /* 0xa4f6 */
            {8'h00}, /* 0xa4f5 */
            {8'h00}, /* 0xa4f4 */
            {8'h00}, /* 0xa4f3 */
            {8'h00}, /* 0xa4f2 */
            {8'h00}, /* 0xa4f1 */
            {8'h00}, /* 0xa4f0 */
            {8'h00}, /* 0xa4ef */
            {8'h00}, /* 0xa4ee */
            {8'h00}, /* 0xa4ed */
            {8'h00}, /* 0xa4ec */
            {8'h00}, /* 0xa4eb */
            {8'h00}, /* 0xa4ea */
            {8'h00}, /* 0xa4e9 */
            {8'h00}, /* 0xa4e8 */
            {8'h00}, /* 0xa4e7 */
            {8'h00}, /* 0xa4e6 */
            {8'h00}, /* 0xa4e5 */
            {8'h00}, /* 0xa4e4 */
            {8'h00}, /* 0xa4e3 */
            {8'h00}, /* 0xa4e2 */
            {8'h00}, /* 0xa4e1 */
            {8'h00}, /* 0xa4e0 */
            {8'h00}, /* 0xa4df */
            {8'h00}, /* 0xa4de */
            {8'h00}, /* 0xa4dd */
            {8'h00}, /* 0xa4dc */
            {8'h00}, /* 0xa4db */
            {8'h00}, /* 0xa4da */
            {8'h00}, /* 0xa4d9 */
            {8'h00}, /* 0xa4d8 */
            {8'h00}, /* 0xa4d7 */
            {8'h00}, /* 0xa4d6 */
            {8'h00}, /* 0xa4d5 */
            {8'h00}, /* 0xa4d4 */
            {8'h00}, /* 0xa4d3 */
            {8'h00}, /* 0xa4d2 */
            {8'h00}, /* 0xa4d1 */
            {8'h00}, /* 0xa4d0 */
            {8'h00}, /* 0xa4cf */
            {8'h00}, /* 0xa4ce */
            {8'h00}, /* 0xa4cd */
            {8'h00}, /* 0xa4cc */
            {8'h00}, /* 0xa4cb */
            {8'h00}, /* 0xa4ca */
            {8'h00}, /* 0xa4c9 */
            {8'h00}, /* 0xa4c8 */
            {8'h00}, /* 0xa4c7 */
            {8'h00}, /* 0xa4c6 */
            {8'h00}, /* 0xa4c5 */
            {8'h00}, /* 0xa4c4 */
            {8'h00}, /* 0xa4c3 */
            {8'h00}, /* 0xa4c2 */
            {8'h00}, /* 0xa4c1 */
            {8'h00}, /* 0xa4c0 */
            {8'h00}, /* 0xa4bf */
            {8'h00}, /* 0xa4be */
            {8'h00}, /* 0xa4bd */
            {8'h00}, /* 0xa4bc */
            {8'h00}, /* 0xa4bb */
            {8'h00}, /* 0xa4ba */
            {8'h00}, /* 0xa4b9 */
            {8'h00}, /* 0xa4b8 */
            {8'h00}, /* 0xa4b7 */
            {8'h00}, /* 0xa4b6 */
            {8'h00}, /* 0xa4b5 */
            {8'h00}, /* 0xa4b4 */
            {8'h00}, /* 0xa4b3 */
            {8'h00}, /* 0xa4b2 */
            {8'h00}, /* 0xa4b1 */
            {8'h00}, /* 0xa4b0 */
            {8'h00}, /* 0xa4af */
            {8'h00}, /* 0xa4ae */
            {8'h00}, /* 0xa4ad */
            {8'h00}, /* 0xa4ac */
            {8'h00}, /* 0xa4ab */
            {8'h00}, /* 0xa4aa */
            {8'h00}, /* 0xa4a9 */
            {8'h00}, /* 0xa4a8 */
            {8'h00}, /* 0xa4a7 */
            {8'h00}, /* 0xa4a6 */
            {8'h00}, /* 0xa4a5 */
            {8'h00}, /* 0xa4a4 */
            {8'h00}, /* 0xa4a3 */
            {8'h00}, /* 0xa4a2 */
            {8'h00}, /* 0xa4a1 */
            {8'h00}, /* 0xa4a0 */
            {8'h00}, /* 0xa49f */
            {8'h00}, /* 0xa49e */
            {8'h00}, /* 0xa49d */
            {8'h00}, /* 0xa49c */
            {8'h00}, /* 0xa49b */
            {8'h00}, /* 0xa49a */
            {8'h00}, /* 0xa499 */
            {8'h00}, /* 0xa498 */
            {8'h00}, /* 0xa497 */
            {8'h00}, /* 0xa496 */
            {8'h00}, /* 0xa495 */
            {8'h00}, /* 0xa494 */
            {8'h00}, /* 0xa493 */
            {8'h00}, /* 0xa492 */
            {8'h00}, /* 0xa491 */
            {8'h00}, /* 0xa490 */
            {8'h00}, /* 0xa48f */
            {8'h00}, /* 0xa48e */
            {8'h00}, /* 0xa48d */
            {8'h00}, /* 0xa48c */
            {8'h00}, /* 0xa48b */
            {8'h00}, /* 0xa48a */
            {8'h00}, /* 0xa489 */
            {8'h00}, /* 0xa488 */
            {8'h00}, /* 0xa487 */
            {8'h00}, /* 0xa486 */
            {8'h00}, /* 0xa485 */
            {8'h00}, /* 0xa484 */
            {8'h00}, /* 0xa483 */
            {8'h00}, /* 0xa482 */
            {8'h00}, /* 0xa481 */
            {8'h00}, /* 0xa480 */
            {8'h00}, /* 0xa47f */
            {8'h00}, /* 0xa47e */
            {8'h00}, /* 0xa47d */
            {8'h00}, /* 0xa47c */
            {8'h00}, /* 0xa47b */
            {8'h00}, /* 0xa47a */
            {8'h00}, /* 0xa479 */
            {8'h00}, /* 0xa478 */
            {8'h00}, /* 0xa477 */
            {8'h00}, /* 0xa476 */
            {8'h00}, /* 0xa475 */
            {8'h00}, /* 0xa474 */
            {8'h00}, /* 0xa473 */
            {8'h00}, /* 0xa472 */
            {8'h00}, /* 0xa471 */
            {8'h00}, /* 0xa470 */
            {8'h00}, /* 0xa46f */
            {8'h00}, /* 0xa46e */
            {8'h00}, /* 0xa46d */
            {8'h00}, /* 0xa46c */
            {8'h00}, /* 0xa46b */
            {8'h00}, /* 0xa46a */
            {8'h00}, /* 0xa469 */
            {8'h00}, /* 0xa468 */
            {8'h00}, /* 0xa467 */
            {8'h00}, /* 0xa466 */
            {8'h00}, /* 0xa465 */
            {8'h00}, /* 0xa464 */
            {8'h00}, /* 0xa463 */
            {8'h00}, /* 0xa462 */
            {8'h00}, /* 0xa461 */
            {8'h00}, /* 0xa460 */
            {8'h00}, /* 0xa45f */
            {8'h00}, /* 0xa45e */
            {8'h00}, /* 0xa45d */
            {8'h00}, /* 0xa45c */
            {8'h00}, /* 0xa45b */
            {8'h00}, /* 0xa45a */
            {8'h00}, /* 0xa459 */
            {8'h00}, /* 0xa458 */
            {8'h00}, /* 0xa457 */
            {8'h00}, /* 0xa456 */
            {8'h00}, /* 0xa455 */
            {8'h00}, /* 0xa454 */
            {8'h00}, /* 0xa453 */
            {8'h00}, /* 0xa452 */
            {8'h00}, /* 0xa451 */
            {8'h00}, /* 0xa450 */
            {8'h00}, /* 0xa44f */
            {8'h00}, /* 0xa44e */
            {8'h00}, /* 0xa44d */
            {8'h00}, /* 0xa44c */
            {8'h00}, /* 0xa44b */
            {8'h00}, /* 0xa44a */
            {8'h00}, /* 0xa449 */
            {8'h00}, /* 0xa448 */
            {8'h00}, /* 0xa447 */
            {8'h00}, /* 0xa446 */
            {8'h00}, /* 0xa445 */
            {8'h00}, /* 0xa444 */
            {8'h00}, /* 0xa443 */
            {8'h00}, /* 0xa442 */
            {8'h00}, /* 0xa441 */
            {8'h00}, /* 0xa440 */
            {8'h00}, /* 0xa43f */
            {8'h00}, /* 0xa43e */
            {8'h00}, /* 0xa43d */
            {8'h00}, /* 0xa43c */
            {8'h00}, /* 0xa43b */
            {8'h00}, /* 0xa43a */
            {8'h00}, /* 0xa439 */
            {8'h00}, /* 0xa438 */
            {8'h00}, /* 0xa437 */
            {8'h00}, /* 0xa436 */
            {8'h00}, /* 0xa435 */
            {8'h00}, /* 0xa434 */
            {8'h00}, /* 0xa433 */
            {8'h00}, /* 0xa432 */
            {8'h00}, /* 0xa431 */
            {8'h00}, /* 0xa430 */
            {8'h00}, /* 0xa42f */
            {8'h00}, /* 0xa42e */
            {8'h00}, /* 0xa42d */
            {8'h00}, /* 0xa42c */
            {8'h00}, /* 0xa42b */
            {8'h00}, /* 0xa42a */
            {8'h00}, /* 0xa429 */
            {8'h00}, /* 0xa428 */
            {8'h00}, /* 0xa427 */
            {8'h00}, /* 0xa426 */
            {8'h00}, /* 0xa425 */
            {8'h00}, /* 0xa424 */
            {8'h00}, /* 0xa423 */
            {8'h00}, /* 0xa422 */
            {8'h00}, /* 0xa421 */
            {8'h00}, /* 0xa420 */
            {8'h00}, /* 0xa41f */
            {8'h00}, /* 0xa41e */
            {8'h00}, /* 0xa41d */
            {8'h00}, /* 0xa41c */
            {8'h00}, /* 0xa41b */
            {8'h00}, /* 0xa41a */
            {8'h00}, /* 0xa419 */
            {8'h00}, /* 0xa418 */
            {8'h00}, /* 0xa417 */
            {8'h00}, /* 0xa416 */
            {8'h00}, /* 0xa415 */
            {8'h00}, /* 0xa414 */
            {8'h00}, /* 0xa413 */
            {8'h00}, /* 0xa412 */
            {8'h00}, /* 0xa411 */
            {8'h00}, /* 0xa410 */
            {8'h00}, /* 0xa40f */
            {8'h00}, /* 0xa40e */
            {8'h00}, /* 0xa40d */
            {8'h00}, /* 0xa40c */
            {8'h00}, /* 0xa40b */
            {8'h00}, /* 0xa40a */
            {8'h00}, /* 0xa409 */
            {8'h00}, /* 0xa408 */
            {8'h00}, /* 0xa407 */
            {8'h00}, /* 0xa406 */
            {8'h00}, /* 0xa405 */
            {8'h00}, /* 0xa404 */
            {8'h00}, /* 0xa403 */
            {8'h00}, /* 0xa402 */
            {8'h00}, /* 0xa401 */
            {8'h00}, /* 0xa400 */
            {8'h00}, /* 0xa3ff */
            {8'h00}, /* 0xa3fe */
            {8'h00}, /* 0xa3fd */
            {8'h00}, /* 0xa3fc */
            {8'h00}, /* 0xa3fb */
            {8'h00}, /* 0xa3fa */
            {8'h00}, /* 0xa3f9 */
            {8'h00}, /* 0xa3f8 */
            {8'h00}, /* 0xa3f7 */
            {8'h00}, /* 0xa3f6 */
            {8'h00}, /* 0xa3f5 */
            {8'h00}, /* 0xa3f4 */
            {8'h00}, /* 0xa3f3 */
            {8'h00}, /* 0xa3f2 */
            {8'h00}, /* 0xa3f1 */
            {8'h00}, /* 0xa3f0 */
            {8'h00}, /* 0xa3ef */
            {8'h00}, /* 0xa3ee */
            {8'h00}, /* 0xa3ed */
            {8'h00}, /* 0xa3ec */
            {8'h00}, /* 0xa3eb */
            {8'h00}, /* 0xa3ea */
            {8'h00}, /* 0xa3e9 */
            {8'h00}, /* 0xa3e8 */
            {8'h00}, /* 0xa3e7 */
            {8'h00}, /* 0xa3e6 */
            {8'h00}, /* 0xa3e5 */
            {8'h00}, /* 0xa3e4 */
            {8'h00}, /* 0xa3e3 */
            {8'h00}, /* 0xa3e2 */
            {8'h00}, /* 0xa3e1 */
            {8'h00}, /* 0xa3e0 */
            {8'h00}, /* 0xa3df */
            {8'h00}, /* 0xa3de */
            {8'h00}, /* 0xa3dd */
            {8'h00}, /* 0xa3dc */
            {8'h00}, /* 0xa3db */
            {8'h00}, /* 0xa3da */
            {8'h00}, /* 0xa3d9 */
            {8'h00}, /* 0xa3d8 */
            {8'h00}, /* 0xa3d7 */
            {8'h00}, /* 0xa3d6 */
            {8'h00}, /* 0xa3d5 */
            {8'h00}, /* 0xa3d4 */
            {8'h00}, /* 0xa3d3 */
            {8'h00}, /* 0xa3d2 */
            {8'h00}, /* 0xa3d1 */
            {8'h00}, /* 0xa3d0 */
            {8'h00}, /* 0xa3cf */
            {8'h00}, /* 0xa3ce */
            {8'h00}, /* 0xa3cd */
            {8'h00}, /* 0xa3cc */
            {8'h00}, /* 0xa3cb */
            {8'h00}, /* 0xa3ca */
            {8'h00}, /* 0xa3c9 */
            {8'h00}, /* 0xa3c8 */
            {8'h00}, /* 0xa3c7 */
            {8'h00}, /* 0xa3c6 */
            {8'h00}, /* 0xa3c5 */
            {8'h00}, /* 0xa3c4 */
            {8'h00}, /* 0xa3c3 */
            {8'h00}, /* 0xa3c2 */
            {8'h00}, /* 0xa3c1 */
            {8'h00}, /* 0xa3c0 */
            {8'h00}, /* 0xa3bf */
            {8'h00}, /* 0xa3be */
            {8'h00}, /* 0xa3bd */
            {8'h00}, /* 0xa3bc */
            {8'h00}, /* 0xa3bb */
            {8'h00}, /* 0xa3ba */
            {8'h00}, /* 0xa3b9 */
            {8'h00}, /* 0xa3b8 */
            {8'h00}, /* 0xa3b7 */
            {8'h00}, /* 0xa3b6 */
            {8'h00}, /* 0xa3b5 */
            {8'h00}, /* 0xa3b4 */
            {8'h00}, /* 0xa3b3 */
            {8'h00}, /* 0xa3b2 */
            {8'h00}, /* 0xa3b1 */
            {8'h00}, /* 0xa3b0 */
            {8'h00}, /* 0xa3af */
            {8'h00}, /* 0xa3ae */
            {8'h00}, /* 0xa3ad */
            {8'h00}, /* 0xa3ac */
            {8'h00}, /* 0xa3ab */
            {8'h00}, /* 0xa3aa */
            {8'h00}, /* 0xa3a9 */
            {8'h00}, /* 0xa3a8 */
            {8'h00}, /* 0xa3a7 */
            {8'h00}, /* 0xa3a6 */
            {8'h00}, /* 0xa3a5 */
            {8'h00}, /* 0xa3a4 */
            {8'h00}, /* 0xa3a3 */
            {8'h00}, /* 0xa3a2 */
            {8'h00}, /* 0xa3a1 */
            {8'h00}, /* 0xa3a0 */
            {8'h00}, /* 0xa39f */
            {8'h00}, /* 0xa39e */
            {8'h00}, /* 0xa39d */
            {8'h00}, /* 0xa39c */
            {8'h00}, /* 0xa39b */
            {8'h00}, /* 0xa39a */
            {8'h00}, /* 0xa399 */
            {8'h00}, /* 0xa398 */
            {8'h00}, /* 0xa397 */
            {8'h00}, /* 0xa396 */
            {8'h00}, /* 0xa395 */
            {8'h00}, /* 0xa394 */
            {8'h00}, /* 0xa393 */
            {8'h00}, /* 0xa392 */
            {8'h00}, /* 0xa391 */
            {8'h00}, /* 0xa390 */
            {8'h00}, /* 0xa38f */
            {8'h00}, /* 0xa38e */
            {8'h00}, /* 0xa38d */
            {8'h00}, /* 0xa38c */
            {8'h00}, /* 0xa38b */
            {8'h00}, /* 0xa38a */
            {8'h00}, /* 0xa389 */
            {8'h00}, /* 0xa388 */
            {8'h00}, /* 0xa387 */
            {8'h00}, /* 0xa386 */
            {8'h00}, /* 0xa385 */
            {8'h00}, /* 0xa384 */
            {8'h00}, /* 0xa383 */
            {8'h00}, /* 0xa382 */
            {8'h00}, /* 0xa381 */
            {8'h00}, /* 0xa380 */
            {8'h00}, /* 0xa37f */
            {8'h00}, /* 0xa37e */
            {8'h00}, /* 0xa37d */
            {8'h00}, /* 0xa37c */
            {8'h00}, /* 0xa37b */
            {8'h00}, /* 0xa37a */
            {8'h00}, /* 0xa379 */
            {8'h00}, /* 0xa378 */
            {8'h00}, /* 0xa377 */
            {8'h00}, /* 0xa376 */
            {8'h00}, /* 0xa375 */
            {8'h00}, /* 0xa374 */
            {8'h00}, /* 0xa373 */
            {8'h00}, /* 0xa372 */
            {8'h00}, /* 0xa371 */
            {8'h00}, /* 0xa370 */
            {8'h00}, /* 0xa36f */
            {8'h00}, /* 0xa36e */
            {8'h00}, /* 0xa36d */
            {8'h00}, /* 0xa36c */
            {8'h00}, /* 0xa36b */
            {8'h00}, /* 0xa36a */
            {8'h00}, /* 0xa369 */
            {8'h00}, /* 0xa368 */
            {8'h00}, /* 0xa367 */
            {8'h00}, /* 0xa366 */
            {8'h00}, /* 0xa365 */
            {8'h00}, /* 0xa364 */
            {8'h00}, /* 0xa363 */
            {8'h00}, /* 0xa362 */
            {8'h00}, /* 0xa361 */
            {8'h00}, /* 0xa360 */
            {8'h00}, /* 0xa35f */
            {8'h00}, /* 0xa35e */
            {8'h00}, /* 0xa35d */
            {8'h00}, /* 0xa35c */
            {8'h00}, /* 0xa35b */
            {8'h00}, /* 0xa35a */
            {8'h00}, /* 0xa359 */
            {8'h00}, /* 0xa358 */
            {8'h00}, /* 0xa357 */
            {8'h00}, /* 0xa356 */
            {8'h00}, /* 0xa355 */
            {8'h00}, /* 0xa354 */
            {8'h00}, /* 0xa353 */
            {8'h00}, /* 0xa352 */
            {8'h00}, /* 0xa351 */
            {8'h00}, /* 0xa350 */
            {8'h00}, /* 0xa34f */
            {8'h00}, /* 0xa34e */
            {8'h00}, /* 0xa34d */
            {8'h00}, /* 0xa34c */
            {8'h00}, /* 0xa34b */
            {8'h00}, /* 0xa34a */
            {8'h00}, /* 0xa349 */
            {8'h00}, /* 0xa348 */
            {8'h00}, /* 0xa347 */
            {8'h00}, /* 0xa346 */
            {8'h00}, /* 0xa345 */
            {8'h00}, /* 0xa344 */
            {8'h00}, /* 0xa343 */
            {8'h00}, /* 0xa342 */
            {8'h00}, /* 0xa341 */
            {8'h00}, /* 0xa340 */
            {8'h00}, /* 0xa33f */
            {8'h00}, /* 0xa33e */
            {8'h00}, /* 0xa33d */
            {8'h00}, /* 0xa33c */
            {8'h00}, /* 0xa33b */
            {8'h00}, /* 0xa33a */
            {8'h00}, /* 0xa339 */
            {8'h00}, /* 0xa338 */
            {8'h00}, /* 0xa337 */
            {8'h00}, /* 0xa336 */
            {8'h00}, /* 0xa335 */
            {8'h00}, /* 0xa334 */
            {8'h00}, /* 0xa333 */
            {8'h00}, /* 0xa332 */
            {8'h00}, /* 0xa331 */
            {8'h00}, /* 0xa330 */
            {8'h00}, /* 0xa32f */
            {8'h00}, /* 0xa32e */
            {8'h00}, /* 0xa32d */
            {8'h00}, /* 0xa32c */
            {8'h00}, /* 0xa32b */
            {8'h00}, /* 0xa32a */
            {8'h00}, /* 0xa329 */
            {8'h00}, /* 0xa328 */
            {8'h00}, /* 0xa327 */
            {8'h00}, /* 0xa326 */
            {8'h00}, /* 0xa325 */
            {8'h00}, /* 0xa324 */
            {8'h00}, /* 0xa323 */
            {8'h00}, /* 0xa322 */
            {8'h00}, /* 0xa321 */
            {8'h00}, /* 0xa320 */
            {8'h00}, /* 0xa31f */
            {8'h00}, /* 0xa31e */
            {8'h00}, /* 0xa31d */
            {8'h00}, /* 0xa31c */
            {8'h00}, /* 0xa31b */
            {8'h00}, /* 0xa31a */
            {8'h00}, /* 0xa319 */
            {8'h00}, /* 0xa318 */
            {8'h00}, /* 0xa317 */
            {8'h00}, /* 0xa316 */
            {8'h00}, /* 0xa315 */
            {8'h00}, /* 0xa314 */
            {8'h00}, /* 0xa313 */
            {8'h00}, /* 0xa312 */
            {8'h00}, /* 0xa311 */
            {8'h00}, /* 0xa310 */
            {8'h00}, /* 0xa30f */
            {8'h00}, /* 0xa30e */
            {8'h00}, /* 0xa30d */
            {8'h00}, /* 0xa30c */
            {8'h00}, /* 0xa30b */
            {8'h00}, /* 0xa30a */
            {8'h00}, /* 0xa309 */
            {8'h00}, /* 0xa308 */
            {8'h00}, /* 0xa307 */
            {8'h00}, /* 0xa306 */
            {8'h00}, /* 0xa305 */
            {8'h00}, /* 0xa304 */
            {8'h00}, /* 0xa303 */
            {8'h00}, /* 0xa302 */
            {8'h00}, /* 0xa301 */
            {8'h00}, /* 0xa300 */
            {8'h00}, /* 0xa2ff */
            {8'h00}, /* 0xa2fe */
            {8'h00}, /* 0xa2fd */
            {8'h00}, /* 0xa2fc */
            {8'h00}, /* 0xa2fb */
            {8'h00}, /* 0xa2fa */
            {8'h00}, /* 0xa2f9 */
            {8'h00}, /* 0xa2f8 */
            {8'h00}, /* 0xa2f7 */
            {8'h00}, /* 0xa2f6 */
            {8'h00}, /* 0xa2f5 */
            {8'h00}, /* 0xa2f4 */
            {8'h00}, /* 0xa2f3 */
            {8'h00}, /* 0xa2f2 */
            {8'h00}, /* 0xa2f1 */
            {8'h00}, /* 0xa2f0 */
            {8'h00}, /* 0xa2ef */
            {8'h00}, /* 0xa2ee */
            {8'h00}, /* 0xa2ed */
            {8'h00}, /* 0xa2ec */
            {8'h00}, /* 0xa2eb */
            {8'h00}, /* 0xa2ea */
            {8'h00}, /* 0xa2e9 */
            {8'h00}, /* 0xa2e8 */
            {8'h00}, /* 0xa2e7 */
            {8'h00}, /* 0xa2e6 */
            {8'h00}, /* 0xa2e5 */
            {8'h00}, /* 0xa2e4 */
            {8'h00}, /* 0xa2e3 */
            {8'h00}, /* 0xa2e2 */
            {8'h00}, /* 0xa2e1 */
            {8'h00}, /* 0xa2e0 */
            {8'h00}, /* 0xa2df */
            {8'h00}, /* 0xa2de */
            {8'h00}, /* 0xa2dd */
            {8'h00}, /* 0xa2dc */
            {8'h00}, /* 0xa2db */
            {8'h00}, /* 0xa2da */
            {8'h00}, /* 0xa2d9 */
            {8'h00}, /* 0xa2d8 */
            {8'h00}, /* 0xa2d7 */
            {8'h00}, /* 0xa2d6 */
            {8'h00}, /* 0xa2d5 */
            {8'h00}, /* 0xa2d4 */
            {8'h00}, /* 0xa2d3 */
            {8'h00}, /* 0xa2d2 */
            {8'h00}, /* 0xa2d1 */
            {8'h00}, /* 0xa2d0 */
            {8'h00}, /* 0xa2cf */
            {8'h00}, /* 0xa2ce */
            {8'h00}, /* 0xa2cd */
            {8'h00}, /* 0xa2cc */
            {8'h00}, /* 0xa2cb */
            {8'h00}, /* 0xa2ca */
            {8'h00}, /* 0xa2c9 */
            {8'h00}, /* 0xa2c8 */
            {8'h00}, /* 0xa2c7 */
            {8'h00}, /* 0xa2c6 */
            {8'h00}, /* 0xa2c5 */
            {8'h00}, /* 0xa2c4 */
            {8'h00}, /* 0xa2c3 */
            {8'h00}, /* 0xa2c2 */
            {8'h00}, /* 0xa2c1 */
            {8'h00}, /* 0xa2c0 */
            {8'h00}, /* 0xa2bf */
            {8'h00}, /* 0xa2be */
            {8'h00}, /* 0xa2bd */
            {8'h00}, /* 0xa2bc */
            {8'h00}, /* 0xa2bb */
            {8'h00}, /* 0xa2ba */
            {8'h00}, /* 0xa2b9 */
            {8'h00}, /* 0xa2b8 */
            {8'h00}, /* 0xa2b7 */
            {8'h00}, /* 0xa2b6 */
            {8'h00}, /* 0xa2b5 */
            {8'h00}, /* 0xa2b4 */
            {8'h00}, /* 0xa2b3 */
            {8'h00}, /* 0xa2b2 */
            {8'h00}, /* 0xa2b1 */
            {8'h00}, /* 0xa2b0 */
            {8'h00}, /* 0xa2af */
            {8'h00}, /* 0xa2ae */
            {8'h00}, /* 0xa2ad */
            {8'h00}, /* 0xa2ac */
            {8'h00}, /* 0xa2ab */
            {8'h00}, /* 0xa2aa */
            {8'h00}, /* 0xa2a9 */
            {8'h00}, /* 0xa2a8 */
            {8'h00}, /* 0xa2a7 */
            {8'h00}, /* 0xa2a6 */
            {8'h00}, /* 0xa2a5 */
            {8'h00}, /* 0xa2a4 */
            {8'h00}, /* 0xa2a3 */
            {8'h00}, /* 0xa2a2 */
            {8'h00}, /* 0xa2a1 */
            {8'h00}, /* 0xa2a0 */
            {8'h00}, /* 0xa29f */
            {8'h00}, /* 0xa29e */
            {8'h00}, /* 0xa29d */
            {8'h00}, /* 0xa29c */
            {8'h00}, /* 0xa29b */
            {8'h00}, /* 0xa29a */
            {8'h00}, /* 0xa299 */
            {8'h00}, /* 0xa298 */
            {8'h00}, /* 0xa297 */
            {8'h00}, /* 0xa296 */
            {8'h00}, /* 0xa295 */
            {8'h00}, /* 0xa294 */
            {8'h00}, /* 0xa293 */
            {8'h00}, /* 0xa292 */
            {8'h00}, /* 0xa291 */
            {8'h00}, /* 0xa290 */
            {8'h00}, /* 0xa28f */
            {8'h00}, /* 0xa28e */
            {8'h00}, /* 0xa28d */
            {8'h00}, /* 0xa28c */
            {8'h00}, /* 0xa28b */
            {8'h00}, /* 0xa28a */
            {8'h00}, /* 0xa289 */
            {8'h00}, /* 0xa288 */
            {8'h00}, /* 0xa287 */
            {8'h00}, /* 0xa286 */
            {8'h00}, /* 0xa285 */
            {8'h00}, /* 0xa284 */
            {8'h00}, /* 0xa283 */
            {8'h00}, /* 0xa282 */
            {8'h00}, /* 0xa281 */
            {8'h00}, /* 0xa280 */
            {8'h00}, /* 0xa27f */
            {8'h00}, /* 0xa27e */
            {8'h00}, /* 0xa27d */
            {8'h00}, /* 0xa27c */
            {8'h00}, /* 0xa27b */
            {8'h00}, /* 0xa27a */
            {8'h00}, /* 0xa279 */
            {8'h00}, /* 0xa278 */
            {8'h00}, /* 0xa277 */
            {8'h00}, /* 0xa276 */
            {8'h00}, /* 0xa275 */
            {8'h00}, /* 0xa274 */
            {8'h00}, /* 0xa273 */
            {8'h00}, /* 0xa272 */
            {8'h00}, /* 0xa271 */
            {8'h00}, /* 0xa270 */
            {8'h00}, /* 0xa26f */
            {8'h00}, /* 0xa26e */
            {8'h00}, /* 0xa26d */
            {8'h00}, /* 0xa26c */
            {8'h00}, /* 0xa26b */
            {8'h00}, /* 0xa26a */
            {8'h00}, /* 0xa269 */
            {8'h00}, /* 0xa268 */
            {8'h00}, /* 0xa267 */
            {8'h00}, /* 0xa266 */
            {8'h00}, /* 0xa265 */
            {8'h00}, /* 0xa264 */
            {8'h00}, /* 0xa263 */
            {8'h00}, /* 0xa262 */
            {8'h00}, /* 0xa261 */
            {8'h00}, /* 0xa260 */
            {8'h00}, /* 0xa25f */
            {8'h00}, /* 0xa25e */
            {8'h00}, /* 0xa25d */
            {8'h00}, /* 0xa25c */
            {8'h00}, /* 0xa25b */
            {8'h00}, /* 0xa25a */
            {8'h00}, /* 0xa259 */
            {8'h00}, /* 0xa258 */
            {8'h00}, /* 0xa257 */
            {8'h00}, /* 0xa256 */
            {8'h00}, /* 0xa255 */
            {8'h00}, /* 0xa254 */
            {8'h00}, /* 0xa253 */
            {8'h00}, /* 0xa252 */
            {8'h00}, /* 0xa251 */
            {8'h00}, /* 0xa250 */
            {8'h00}, /* 0xa24f */
            {8'h00}, /* 0xa24e */
            {8'h00}, /* 0xa24d */
            {8'h00}, /* 0xa24c */
            {8'h00}, /* 0xa24b */
            {8'h00}, /* 0xa24a */
            {8'h00}, /* 0xa249 */
            {8'h00}, /* 0xa248 */
            {8'h00}, /* 0xa247 */
            {8'h00}, /* 0xa246 */
            {8'h00}, /* 0xa245 */
            {8'h00}, /* 0xa244 */
            {8'h00}, /* 0xa243 */
            {8'h00}, /* 0xa242 */
            {8'h00}, /* 0xa241 */
            {8'h00}, /* 0xa240 */
            {8'h00}, /* 0xa23f */
            {8'h00}, /* 0xa23e */
            {8'h00}, /* 0xa23d */
            {8'h00}, /* 0xa23c */
            {8'h00}, /* 0xa23b */
            {8'h00}, /* 0xa23a */
            {8'h00}, /* 0xa239 */
            {8'h00}, /* 0xa238 */
            {8'h00}, /* 0xa237 */
            {8'h00}, /* 0xa236 */
            {8'h00}, /* 0xa235 */
            {8'h00}, /* 0xa234 */
            {8'h00}, /* 0xa233 */
            {8'h00}, /* 0xa232 */
            {8'h00}, /* 0xa231 */
            {8'h00}, /* 0xa230 */
            {8'h00}, /* 0xa22f */
            {8'h00}, /* 0xa22e */
            {8'h00}, /* 0xa22d */
            {8'h00}, /* 0xa22c */
            {8'h00}, /* 0xa22b */
            {8'h00}, /* 0xa22a */
            {8'h00}, /* 0xa229 */
            {8'h00}, /* 0xa228 */
            {8'h00}, /* 0xa227 */
            {8'h00}, /* 0xa226 */
            {8'h00}, /* 0xa225 */
            {8'h00}, /* 0xa224 */
            {8'h00}, /* 0xa223 */
            {8'h00}, /* 0xa222 */
            {8'h00}, /* 0xa221 */
            {8'h00}, /* 0xa220 */
            {8'h00}, /* 0xa21f */
            {8'h00}, /* 0xa21e */
            {8'h00}, /* 0xa21d */
            {8'h00}, /* 0xa21c */
            {8'h00}, /* 0xa21b */
            {8'h00}, /* 0xa21a */
            {8'h00}, /* 0xa219 */
            {8'h00}, /* 0xa218 */
            {8'h00}, /* 0xa217 */
            {8'h00}, /* 0xa216 */
            {8'h00}, /* 0xa215 */
            {8'h00}, /* 0xa214 */
            {8'h00}, /* 0xa213 */
            {8'h00}, /* 0xa212 */
            {8'h00}, /* 0xa211 */
            {8'h00}, /* 0xa210 */
            {8'h00}, /* 0xa20f */
            {8'h00}, /* 0xa20e */
            {8'h00}, /* 0xa20d */
            {8'h00}, /* 0xa20c */
            {8'h00}, /* 0xa20b */
            {8'h00}, /* 0xa20a */
            {8'h00}, /* 0xa209 */
            {8'h00}, /* 0xa208 */
            {8'h00}, /* 0xa207 */
            {8'h00}, /* 0xa206 */
            {8'h00}, /* 0xa205 */
            {8'h00}, /* 0xa204 */
            {8'h00}, /* 0xa203 */
            {8'h00}, /* 0xa202 */
            {8'h00}, /* 0xa201 */
            {8'h00}, /* 0xa200 */
            {8'h00}, /* 0xa1ff */
            {8'h00}, /* 0xa1fe */
            {8'h00}, /* 0xa1fd */
            {8'h00}, /* 0xa1fc */
            {8'h00}, /* 0xa1fb */
            {8'h00}, /* 0xa1fa */
            {8'h00}, /* 0xa1f9 */
            {8'h00}, /* 0xa1f8 */
            {8'h00}, /* 0xa1f7 */
            {8'h00}, /* 0xa1f6 */
            {8'h00}, /* 0xa1f5 */
            {8'h00}, /* 0xa1f4 */
            {8'h00}, /* 0xa1f3 */
            {8'h00}, /* 0xa1f2 */
            {8'h00}, /* 0xa1f1 */
            {8'h00}, /* 0xa1f0 */
            {8'h00}, /* 0xa1ef */
            {8'h00}, /* 0xa1ee */
            {8'h00}, /* 0xa1ed */
            {8'h00}, /* 0xa1ec */
            {8'h00}, /* 0xa1eb */
            {8'h00}, /* 0xa1ea */
            {8'h00}, /* 0xa1e9 */
            {8'h00}, /* 0xa1e8 */
            {8'h00}, /* 0xa1e7 */
            {8'h00}, /* 0xa1e6 */
            {8'h00}, /* 0xa1e5 */
            {8'h00}, /* 0xa1e4 */
            {8'h00}, /* 0xa1e3 */
            {8'h00}, /* 0xa1e2 */
            {8'h00}, /* 0xa1e1 */
            {8'h00}, /* 0xa1e0 */
            {8'h00}, /* 0xa1df */
            {8'h00}, /* 0xa1de */
            {8'h00}, /* 0xa1dd */
            {8'h00}, /* 0xa1dc */
            {8'h00}, /* 0xa1db */
            {8'h00}, /* 0xa1da */
            {8'h00}, /* 0xa1d9 */
            {8'h00}, /* 0xa1d8 */
            {8'h00}, /* 0xa1d7 */
            {8'h00}, /* 0xa1d6 */
            {8'h00}, /* 0xa1d5 */
            {8'h00}, /* 0xa1d4 */
            {8'h00}, /* 0xa1d3 */
            {8'h00}, /* 0xa1d2 */
            {8'h00}, /* 0xa1d1 */
            {8'h00}, /* 0xa1d0 */
            {8'h00}, /* 0xa1cf */
            {8'h00}, /* 0xa1ce */
            {8'h00}, /* 0xa1cd */
            {8'h00}, /* 0xa1cc */
            {8'h00}, /* 0xa1cb */
            {8'h00}, /* 0xa1ca */
            {8'h00}, /* 0xa1c9 */
            {8'h00}, /* 0xa1c8 */
            {8'h00}, /* 0xa1c7 */
            {8'h00}, /* 0xa1c6 */
            {8'h00}, /* 0xa1c5 */
            {8'h00}, /* 0xa1c4 */
            {8'h00}, /* 0xa1c3 */
            {8'h00}, /* 0xa1c2 */
            {8'h00}, /* 0xa1c1 */
            {8'h00}, /* 0xa1c0 */
            {8'h00}, /* 0xa1bf */
            {8'h00}, /* 0xa1be */
            {8'h00}, /* 0xa1bd */
            {8'h00}, /* 0xa1bc */
            {8'h00}, /* 0xa1bb */
            {8'h00}, /* 0xa1ba */
            {8'h00}, /* 0xa1b9 */
            {8'h00}, /* 0xa1b8 */
            {8'h00}, /* 0xa1b7 */
            {8'h00}, /* 0xa1b6 */
            {8'h00}, /* 0xa1b5 */
            {8'h00}, /* 0xa1b4 */
            {8'h00}, /* 0xa1b3 */
            {8'h00}, /* 0xa1b2 */
            {8'h00}, /* 0xa1b1 */
            {8'h00}, /* 0xa1b0 */
            {8'h00}, /* 0xa1af */
            {8'h00}, /* 0xa1ae */
            {8'h00}, /* 0xa1ad */
            {8'h00}, /* 0xa1ac */
            {8'h00}, /* 0xa1ab */
            {8'h00}, /* 0xa1aa */
            {8'h00}, /* 0xa1a9 */
            {8'h00}, /* 0xa1a8 */
            {8'h00}, /* 0xa1a7 */
            {8'h00}, /* 0xa1a6 */
            {8'h00}, /* 0xa1a5 */
            {8'h00}, /* 0xa1a4 */
            {8'h00}, /* 0xa1a3 */
            {8'h00}, /* 0xa1a2 */
            {8'h00}, /* 0xa1a1 */
            {8'h00}, /* 0xa1a0 */
            {8'h00}, /* 0xa19f */
            {8'h00}, /* 0xa19e */
            {8'h00}, /* 0xa19d */
            {8'h00}, /* 0xa19c */
            {8'h00}, /* 0xa19b */
            {8'h00}, /* 0xa19a */
            {8'h00}, /* 0xa199 */
            {8'h00}, /* 0xa198 */
            {8'h00}, /* 0xa197 */
            {8'h00}, /* 0xa196 */
            {8'h00}, /* 0xa195 */
            {8'h00}, /* 0xa194 */
            {8'h00}, /* 0xa193 */
            {8'h00}, /* 0xa192 */
            {8'h00}, /* 0xa191 */
            {8'h00}, /* 0xa190 */
            {8'h00}, /* 0xa18f */
            {8'h00}, /* 0xa18e */
            {8'h00}, /* 0xa18d */
            {8'h00}, /* 0xa18c */
            {8'h00}, /* 0xa18b */
            {8'h00}, /* 0xa18a */
            {8'h00}, /* 0xa189 */
            {8'h00}, /* 0xa188 */
            {8'h00}, /* 0xa187 */
            {8'h00}, /* 0xa186 */
            {8'h00}, /* 0xa185 */
            {8'h00}, /* 0xa184 */
            {8'h00}, /* 0xa183 */
            {8'h00}, /* 0xa182 */
            {8'h00}, /* 0xa181 */
            {8'h00}, /* 0xa180 */
            {8'h00}, /* 0xa17f */
            {8'h00}, /* 0xa17e */
            {8'h00}, /* 0xa17d */
            {8'h00}, /* 0xa17c */
            {8'h00}, /* 0xa17b */
            {8'h00}, /* 0xa17a */
            {8'h00}, /* 0xa179 */
            {8'h00}, /* 0xa178 */
            {8'h00}, /* 0xa177 */
            {8'h00}, /* 0xa176 */
            {8'h00}, /* 0xa175 */
            {8'h00}, /* 0xa174 */
            {8'h00}, /* 0xa173 */
            {8'h00}, /* 0xa172 */
            {8'h00}, /* 0xa171 */
            {8'h00}, /* 0xa170 */
            {8'h00}, /* 0xa16f */
            {8'h00}, /* 0xa16e */
            {8'h00}, /* 0xa16d */
            {8'h00}, /* 0xa16c */
            {8'h00}, /* 0xa16b */
            {8'h00}, /* 0xa16a */
            {8'h00}, /* 0xa169 */
            {8'h00}, /* 0xa168 */
            {8'h00}, /* 0xa167 */
            {8'h00}, /* 0xa166 */
            {8'h00}, /* 0xa165 */
            {8'h00}, /* 0xa164 */
            {8'h00}, /* 0xa163 */
            {8'h00}, /* 0xa162 */
            {8'h00}, /* 0xa161 */
            {8'h00}, /* 0xa160 */
            {8'h00}, /* 0xa15f */
            {8'h00}, /* 0xa15e */
            {8'h00}, /* 0xa15d */
            {8'h00}, /* 0xa15c */
            {8'h00}, /* 0xa15b */
            {8'h00}, /* 0xa15a */
            {8'h00}, /* 0xa159 */
            {8'h00}, /* 0xa158 */
            {8'h00}, /* 0xa157 */
            {8'h00}, /* 0xa156 */
            {8'h00}, /* 0xa155 */
            {8'h00}, /* 0xa154 */
            {8'h00}, /* 0xa153 */
            {8'h00}, /* 0xa152 */
            {8'h00}, /* 0xa151 */
            {8'h00}, /* 0xa150 */
            {8'h00}, /* 0xa14f */
            {8'h00}, /* 0xa14e */
            {8'h00}, /* 0xa14d */
            {8'h00}, /* 0xa14c */
            {8'h00}, /* 0xa14b */
            {8'h00}, /* 0xa14a */
            {8'h00}, /* 0xa149 */
            {8'h00}, /* 0xa148 */
            {8'h00}, /* 0xa147 */
            {8'h00}, /* 0xa146 */
            {8'h00}, /* 0xa145 */
            {8'h00}, /* 0xa144 */
            {8'h00}, /* 0xa143 */
            {8'h00}, /* 0xa142 */
            {8'h00}, /* 0xa141 */
            {8'h00}, /* 0xa140 */
            {8'h00}, /* 0xa13f */
            {8'h00}, /* 0xa13e */
            {8'h00}, /* 0xa13d */
            {8'h00}, /* 0xa13c */
            {8'h00}, /* 0xa13b */
            {8'h00}, /* 0xa13a */
            {8'h00}, /* 0xa139 */
            {8'h00}, /* 0xa138 */
            {8'h00}, /* 0xa137 */
            {8'h00}, /* 0xa136 */
            {8'h00}, /* 0xa135 */
            {8'h00}, /* 0xa134 */
            {8'h00}, /* 0xa133 */
            {8'h00}, /* 0xa132 */
            {8'h00}, /* 0xa131 */
            {8'h00}, /* 0xa130 */
            {8'h00}, /* 0xa12f */
            {8'h00}, /* 0xa12e */
            {8'h00}, /* 0xa12d */
            {8'h00}, /* 0xa12c */
            {8'h00}, /* 0xa12b */
            {8'h00}, /* 0xa12a */
            {8'h00}, /* 0xa129 */
            {8'h00}, /* 0xa128 */
            {8'h00}, /* 0xa127 */
            {8'h00}, /* 0xa126 */
            {8'h00}, /* 0xa125 */
            {8'h00}, /* 0xa124 */
            {8'h00}, /* 0xa123 */
            {8'h00}, /* 0xa122 */
            {8'h00}, /* 0xa121 */
            {8'h00}, /* 0xa120 */
            {8'h00}, /* 0xa11f */
            {8'h00}, /* 0xa11e */
            {8'h00}, /* 0xa11d */
            {8'h00}, /* 0xa11c */
            {8'h00}, /* 0xa11b */
            {8'h00}, /* 0xa11a */
            {8'h00}, /* 0xa119 */
            {8'h00}, /* 0xa118 */
            {8'h00}, /* 0xa117 */
            {8'h00}, /* 0xa116 */
            {8'h00}, /* 0xa115 */
            {8'h00}, /* 0xa114 */
            {8'h00}, /* 0xa113 */
            {8'h00}, /* 0xa112 */
            {8'h00}, /* 0xa111 */
            {8'h00}, /* 0xa110 */
            {8'h00}, /* 0xa10f */
            {8'h00}, /* 0xa10e */
            {8'h00}, /* 0xa10d */
            {8'h00}, /* 0xa10c */
            {8'h00}, /* 0xa10b */
            {8'h00}, /* 0xa10a */
            {8'h00}, /* 0xa109 */
            {8'h00}, /* 0xa108 */
            {8'h00}, /* 0xa107 */
            {8'h00}, /* 0xa106 */
            {8'h00}, /* 0xa105 */
            {8'h00}, /* 0xa104 */
            {8'h00}, /* 0xa103 */
            {8'h00}, /* 0xa102 */
            {8'h00}, /* 0xa101 */
            {8'h00}, /* 0xa100 */
            {8'h00}, /* 0xa0ff */
            {8'h00}, /* 0xa0fe */
            {8'h00}, /* 0xa0fd */
            {8'h00}, /* 0xa0fc */
            {8'h00}, /* 0xa0fb */
            {8'h00}, /* 0xa0fa */
            {8'h00}, /* 0xa0f9 */
            {8'h00}, /* 0xa0f8 */
            {8'h00}, /* 0xa0f7 */
            {8'h00}, /* 0xa0f6 */
            {8'h00}, /* 0xa0f5 */
            {8'h00}, /* 0xa0f4 */
            {8'h00}, /* 0xa0f3 */
            {8'h00}, /* 0xa0f2 */
            {8'h00}, /* 0xa0f1 */
            {8'h00}, /* 0xa0f0 */
            {8'h00}, /* 0xa0ef */
            {8'h00}, /* 0xa0ee */
            {8'h00}, /* 0xa0ed */
            {8'h00}, /* 0xa0ec */
            {8'h00}, /* 0xa0eb */
            {8'h00}, /* 0xa0ea */
            {8'h00}, /* 0xa0e9 */
            {8'h00}, /* 0xa0e8 */
            {8'h00}, /* 0xa0e7 */
            {8'h00}, /* 0xa0e6 */
            {8'h00}, /* 0xa0e5 */
            {8'h00}, /* 0xa0e4 */
            {8'h00}, /* 0xa0e3 */
            {8'h00}, /* 0xa0e2 */
            {8'h00}, /* 0xa0e1 */
            {8'h00}, /* 0xa0e0 */
            {8'h00}, /* 0xa0df */
            {8'h00}, /* 0xa0de */
            {8'h00}, /* 0xa0dd */
            {8'h00}, /* 0xa0dc */
            {8'h00}, /* 0xa0db */
            {8'h00}, /* 0xa0da */
            {8'h00}, /* 0xa0d9 */
            {8'h00}, /* 0xa0d8 */
            {8'h00}, /* 0xa0d7 */
            {8'h00}, /* 0xa0d6 */
            {8'h00}, /* 0xa0d5 */
            {8'h00}, /* 0xa0d4 */
            {8'h00}, /* 0xa0d3 */
            {8'h00}, /* 0xa0d2 */
            {8'h00}, /* 0xa0d1 */
            {8'h00}, /* 0xa0d0 */
            {8'h00}, /* 0xa0cf */
            {8'h00}, /* 0xa0ce */
            {8'h00}, /* 0xa0cd */
            {8'h00}, /* 0xa0cc */
            {8'h00}, /* 0xa0cb */
            {8'h00}, /* 0xa0ca */
            {8'h00}, /* 0xa0c9 */
            {8'h00}, /* 0xa0c8 */
            {8'h00}, /* 0xa0c7 */
            {8'h00}, /* 0xa0c6 */
            {8'h00}, /* 0xa0c5 */
            {8'h00}, /* 0xa0c4 */
            {8'h00}, /* 0xa0c3 */
            {8'h00}, /* 0xa0c2 */
            {8'h00}, /* 0xa0c1 */
            {8'h00}, /* 0xa0c0 */
            {8'h00}, /* 0xa0bf */
            {8'h00}, /* 0xa0be */
            {8'h00}, /* 0xa0bd */
            {8'h00}, /* 0xa0bc */
            {8'h00}, /* 0xa0bb */
            {8'h00}, /* 0xa0ba */
            {8'h00}, /* 0xa0b9 */
            {8'h00}, /* 0xa0b8 */
            {8'h00}, /* 0xa0b7 */
            {8'h00}, /* 0xa0b6 */
            {8'h00}, /* 0xa0b5 */
            {8'h00}, /* 0xa0b4 */
            {8'h00}, /* 0xa0b3 */
            {8'h00}, /* 0xa0b2 */
            {8'h00}, /* 0xa0b1 */
            {8'h00}, /* 0xa0b0 */
            {8'h00}, /* 0xa0af */
            {8'h00}, /* 0xa0ae */
            {8'h00}, /* 0xa0ad */
            {8'h00}, /* 0xa0ac */
            {8'h00}, /* 0xa0ab */
            {8'h00}, /* 0xa0aa */
            {8'h00}, /* 0xa0a9 */
            {8'h00}, /* 0xa0a8 */
            {8'h00}, /* 0xa0a7 */
            {8'h00}, /* 0xa0a6 */
            {8'h00}, /* 0xa0a5 */
            {8'h00}, /* 0xa0a4 */
            {8'h00}, /* 0xa0a3 */
            {8'h00}, /* 0xa0a2 */
            {8'h00}, /* 0xa0a1 */
            {8'h00}, /* 0xa0a0 */
            {8'h00}, /* 0xa09f */
            {8'h00}, /* 0xa09e */
            {8'h00}, /* 0xa09d */
            {8'h00}, /* 0xa09c */
            {8'h00}, /* 0xa09b */
            {8'h00}, /* 0xa09a */
            {8'h00}, /* 0xa099 */
            {8'h00}, /* 0xa098 */
            {8'h00}, /* 0xa097 */
            {8'h00}, /* 0xa096 */
            {8'h00}, /* 0xa095 */
            {8'h00}, /* 0xa094 */
            {8'h00}, /* 0xa093 */
            {8'h00}, /* 0xa092 */
            {8'h00}, /* 0xa091 */
            {8'h00}, /* 0xa090 */
            {8'h00}, /* 0xa08f */
            {8'h00}, /* 0xa08e */
            {8'h00}, /* 0xa08d */
            {8'h00}, /* 0xa08c */
            {8'h00}, /* 0xa08b */
            {8'h00}, /* 0xa08a */
            {8'h00}, /* 0xa089 */
            {8'h00}, /* 0xa088 */
            {8'h00}, /* 0xa087 */
            {8'h00}, /* 0xa086 */
            {8'h00}, /* 0xa085 */
            {8'h00}, /* 0xa084 */
            {8'h00}, /* 0xa083 */
            {8'h00}, /* 0xa082 */
            {8'h00}, /* 0xa081 */
            {8'h00}, /* 0xa080 */
            {8'h00}, /* 0xa07f */
            {8'h00}, /* 0xa07e */
            {8'h00}, /* 0xa07d */
            {8'h00}, /* 0xa07c */
            {8'h00}, /* 0xa07b */
            {8'h00}, /* 0xa07a */
            {8'h00}, /* 0xa079 */
            {8'h00}, /* 0xa078 */
            {8'h00}, /* 0xa077 */
            {8'h00}, /* 0xa076 */
            {8'h00}, /* 0xa075 */
            {8'h00}, /* 0xa074 */
            {8'h00}, /* 0xa073 */
            {8'h00}, /* 0xa072 */
            {8'h00}, /* 0xa071 */
            {8'h00}, /* 0xa070 */
            {8'h00}, /* 0xa06f */
            {8'h00}, /* 0xa06e */
            {8'h00}, /* 0xa06d */
            {8'h00}, /* 0xa06c */
            {8'h00}, /* 0xa06b */
            {8'h00}, /* 0xa06a */
            {8'h00}, /* 0xa069 */
            {8'h00}, /* 0xa068 */
            {8'h00}, /* 0xa067 */
            {8'h00}, /* 0xa066 */
            {8'h00}, /* 0xa065 */
            {8'h00}, /* 0xa064 */
            {8'h00}, /* 0xa063 */
            {8'h00}, /* 0xa062 */
            {8'h00}, /* 0xa061 */
            {8'h00}, /* 0xa060 */
            {8'h00}, /* 0xa05f */
            {8'h00}, /* 0xa05e */
            {8'h00}, /* 0xa05d */
            {8'h00}, /* 0xa05c */
            {8'h00}, /* 0xa05b */
            {8'h00}, /* 0xa05a */
            {8'h00}, /* 0xa059 */
            {8'h00}, /* 0xa058 */
            {8'h00}, /* 0xa057 */
            {8'h00}, /* 0xa056 */
            {8'h00}, /* 0xa055 */
            {8'h00}, /* 0xa054 */
            {8'h00}, /* 0xa053 */
            {8'h00}, /* 0xa052 */
            {8'h00}, /* 0xa051 */
            {8'h00}, /* 0xa050 */
            {8'h00}, /* 0xa04f */
            {8'h00}, /* 0xa04e */
            {8'h00}, /* 0xa04d */
            {8'h00}, /* 0xa04c */
            {8'h00}, /* 0xa04b */
            {8'h00}, /* 0xa04a */
            {8'h00}, /* 0xa049 */
            {8'h00}, /* 0xa048 */
            {8'h00}, /* 0xa047 */
            {8'h00}, /* 0xa046 */
            {8'h00}, /* 0xa045 */
            {8'h00}, /* 0xa044 */
            {8'h00}, /* 0xa043 */
            {8'h00}, /* 0xa042 */
            {8'h00}, /* 0xa041 */
            {8'h00}, /* 0xa040 */
            {8'h00}, /* 0xa03f */
            {8'h00}, /* 0xa03e */
            {8'h00}, /* 0xa03d */
            {8'h00}, /* 0xa03c */
            {8'h00}, /* 0xa03b */
            {8'h00}, /* 0xa03a */
            {8'h00}, /* 0xa039 */
            {8'h00}, /* 0xa038 */
            {8'h00}, /* 0xa037 */
            {8'h00}, /* 0xa036 */
            {8'h00}, /* 0xa035 */
            {8'h00}, /* 0xa034 */
            {8'h00}, /* 0xa033 */
            {8'h00}, /* 0xa032 */
            {8'h00}, /* 0xa031 */
            {8'h00}, /* 0xa030 */
            {8'h00}, /* 0xa02f */
            {8'h00}, /* 0xa02e */
            {8'h00}, /* 0xa02d */
            {8'h00}, /* 0xa02c */
            {8'h00}, /* 0xa02b */
            {8'h00}, /* 0xa02a */
            {8'h00}, /* 0xa029 */
            {8'h00}, /* 0xa028 */
            {8'h00}, /* 0xa027 */
            {8'h00}, /* 0xa026 */
            {8'h00}, /* 0xa025 */
            {8'h00}, /* 0xa024 */
            {8'h00}, /* 0xa023 */
            {8'h00}, /* 0xa022 */
            {8'h00}, /* 0xa021 */
            {8'h00}, /* 0xa020 */
            {8'h00}, /* 0xa01f */
            {8'h00}, /* 0xa01e */
            {8'h00}, /* 0xa01d */
            {8'h00}, /* 0xa01c */
            {8'h00}, /* 0xa01b */
            {8'h00}, /* 0xa01a */
            {8'h00}, /* 0xa019 */
            {8'h00}, /* 0xa018 */
            {8'h00}, /* 0xa017 */
            {8'h00}, /* 0xa016 */
            {8'h00}, /* 0xa015 */
            {8'h00}, /* 0xa014 */
            {8'h00}, /* 0xa013 */
            {8'h00}, /* 0xa012 */
            {8'h00}, /* 0xa011 */
            {8'h00}, /* 0xa010 */
            {8'h00}, /* 0xa00f */
            {8'h00}, /* 0xa00e */
            {8'h00}, /* 0xa00d */
            {8'h00}, /* 0xa00c */
            {8'h00}, /* 0xa00b */
            {8'h00}, /* 0xa00a */
            {8'h00}, /* 0xa009 */
            {8'h00}, /* 0xa008 */
            {8'h00}, /* 0xa007 */
            {8'h00}, /* 0xa006 */
            {8'h00}, /* 0xa005 */
            {8'h00}, /* 0xa004 */
            {8'h00}, /* 0xa003 */
            {8'h00}, /* 0xa002 */
            {8'h00}, /* 0xa001 */
            {8'h00}, /* 0xa000 */
            {8'h00}, /* 0x9fff */
            {8'h00}, /* 0x9ffe */
            {8'h00}, /* 0x9ffd */
            {8'h00}, /* 0x9ffc */
            {8'h00}, /* 0x9ffb */
            {8'h00}, /* 0x9ffa */
            {8'h00}, /* 0x9ff9 */
            {8'h00}, /* 0x9ff8 */
            {8'h00}, /* 0x9ff7 */
            {8'h00}, /* 0x9ff6 */
            {8'h00}, /* 0x9ff5 */
            {8'h00}, /* 0x9ff4 */
            {8'h00}, /* 0x9ff3 */
            {8'h00}, /* 0x9ff2 */
            {8'h00}, /* 0x9ff1 */
            {8'h00}, /* 0x9ff0 */
            {8'h00}, /* 0x9fef */
            {8'h00}, /* 0x9fee */
            {8'h00}, /* 0x9fed */
            {8'h00}, /* 0x9fec */
            {8'h00}, /* 0x9feb */
            {8'h00}, /* 0x9fea */
            {8'h00}, /* 0x9fe9 */
            {8'h00}, /* 0x9fe8 */
            {8'h00}, /* 0x9fe7 */
            {8'h00}, /* 0x9fe6 */
            {8'h00}, /* 0x9fe5 */
            {8'h00}, /* 0x9fe4 */
            {8'h00}, /* 0x9fe3 */
            {8'h00}, /* 0x9fe2 */
            {8'h00}, /* 0x9fe1 */
            {8'h00}, /* 0x9fe0 */
            {8'h00}, /* 0x9fdf */
            {8'h00}, /* 0x9fde */
            {8'h00}, /* 0x9fdd */
            {8'h00}, /* 0x9fdc */
            {8'h00}, /* 0x9fdb */
            {8'h00}, /* 0x9fda */
            {8'h00}, /* 0x9fd9 */
            {8'h00}, /* 0x9fd8 */
            {8'h00}, /* 0x9fd7 */
            {8'h00}, /* 0x9fd6 */
            {8'h00}, /* 0x9fd5 */
            {8'h00}, /* 0x9fd4 */
            {8'h00}, /* 0x9fd3 */
            {8'h00}, /* 0x9fd2 */
            {8'h00}, /* 0x9fd1 */
            {8'h00}, /* 0x9fd0 */
            {8'h00}, /* 0x9fcf */
            {8'h00}, /* 0x9fce */
            {8'h00}, /* 0x9fcd */
            {8'h00}, /* 0x9fcc */
            {8'h00}, /* 0x9fcb */
            {8'h00}, /* 0x9fca */
            {8'h00}, /* 0x9fc9 */
            {8'h00}, /* 0x9fc8 */
            {8'h00}, /* 0x9fc7 */
            {8'h00}, /* 0x9fc6 */
            {8'h00}, /* 0x9fc5 */
            {8'h00}, /* 0x9fc4 */
            {8'h00}, /* 0x9fc3 */
            {8'h00}, /* 0x9fc2 */
            {8'h00}, /* 0x9fc1 */
            {8'h00}, /* 0x9fc0 */
            {8'h00}, /* 0x9fbf */
            {8'h00}, /* 0x9fbe */
            {8'h00}, /* 0x9fbd */
            {8'h00}, /* 0x9fbc */
            {8'h00}, /* 0x9fbb */
            {8'h00}, /* 0x9fba */
            {8'h00}, /* 0x9fb9 */
            {8'h00}, /* 0x9fb8 */
            {8'h00}, /* 0x9fb7 */
            {8'h00}, /* 0x9fb6 */
            {8'h00}, /* 0x9fb5 */
            {8'h00}, /* 0x9fb4 */
            {8'h00}, /* 0x9fb3 */
            {8'h00}, /* 0x9fb2 */
            {8'h00}, /* 0x9fb1 */
            {8'h00}, /* 0x9fb0 */
            {8'h00}, /* 0x9faf */
            {8'h00}, /* 0x9fae */
            {8'h00}, /* 0x9fad */
            {8'h00}, /* 0x9fac */
            {8'h00}, /* 0x9fab */
            {8'h00}, /* 0x9faa */
            {8'h00}, /* 0x9fa9 */
            {8'h00}, /* 0x9fa8 */
            {8'h00}, /* 0x9fa7 */
            {8'h00}, /* 0x9fa6 */
            {8'h00}, /* 0x9fa5 */
            {8'h00}, /* 0x9fa4 */
            {8'h00}, /* 0x9fa3 */
            {8'h00}, /* 0x9fa2 */
            {8'h00}, /* 0x9fa1 */
            {8'h00}, /* 0x9fa0 */
            {8'h00}, /* 0x9f9f */
            {8'h00}, /* 0x9f9e */
            {8'h00}, /* 0x9f9d */
            {8'h00}, /* 0x9f9c */
            {8'h00}, /* 0x9f9b */
            {8'h00}, /* 0x9f9a */
            {8'h00}, /* 0x9f99 */
            {8'h00}, /* 0x9f98 */
            {8'h00}, /* 0x9f97 */
            {8'h00}, /* 0x9f96 */
            {8'h00}, /* 0x9f95 */
            {8'h00}, /* 0x9f94 */
            {8'h00}, /* 0x9f93 */
            {8'h00}, /* 0x9f92 */
            {8'h00}, /* 0x9f91 */
            {8'h00}, /* 0x9f90 */
            {8'h00}, /* 0x9f8f */
            {8'h00}, /* 0x9f8e */
            {8'h00}, /* 0x9f8d */
            {8'h00}, /* 0x9f8c */
            {8'h00}, /* 0x9f8b */
            {8'h00}, /* 0x9f8a */
            {8'h00}, /* 0x9f89 */
            {8'h00}, /* 0x9f88 */
            {8'h00}, /* 0x9f87 */
            {8'h00}, /* 0x9f86 */
            {8'h00}, /* 0x9f85 */
            {8'h00}, /* 0x9f84 */
            {8'h00}, /* 0x9f83 */
            {8'h00}, /* 0x9f82 */
            {8'h00}, /* 0x9f81 */
            {8'h00}, /* 0x9f80 */
            {8'h00}, /* 0x9f7f */
            {8'h00}, /* 0x9f7e */
            {8'h00}, /* 0x9f7d */
            {8'h00}, /* 0x9f7c */
            {8'h00}, /* 0x9f7b */
            {8'h00}, /* 0x9f7a */
            {8'h00}, /* 0x9f79 */
            {8'h00}, /* 0x9f78 */
            {8'h00}, /* 0x9f77 */
            {8'h00}, /* 0x9f76 */
            {8'h00}, /* 0x9f75 */
            {8'h00}, /* 0x9f74 */
            {8'h00}, /* 0x9f73 */
            {8'h00}, /* 0x9f72 */
            {8'h00}, /* 0x9f71 */
            {8'h00}, /* 0x9f70 */
            {8'h00}, /* 0x9f6f */
            {8'h00}, /* 0x9f6e */
            {8'h00}, /* 0x9f6d */
            {8'h00}, /* 0x9f6c */
            {8'h00}, /* 0x9f6b */
            {8'h00}, /* 0x9f6a */
            {8'h00}, /* 0x9f69 */
            {8'h00}, /* 0x9f68 */
            {8'h00}, /* 0x9f67 */
            {8'h00}, /* 0x9f66 */
            {8'h00}, /* 0x9f65 */
            {8'h00}, /* 0x9f64 */
            {8'h00}, /* 0x9f63 */
            {8'h00}, /* 0x9f62 */
            {8'h00}, /* 0x9f61 */
            {8'h00}, /* 0x9f60 */
            {8'h00}, /* 0x9f5f */
            {8'h00}, /* 0x9f5e */
            {8'h00}, /* 0x9f5d */
            {8'h00}, /* 0x9f5c */
            {8'h00}, /* 0x9f5b */
            {8'h00}, /* 0x9f5a */
            {8'h00}, /* 0x9f59 */
            {8'h00}, /* 0x9f58 */
            {8'h00}, /* 0x9f57 */
            {8'h00}, /* 0x9f56 */
            {8'h00}, /* 0x9f55 */
            {8'h00}, /* 0x9f54 */
            {8'h00}, /* 0x9f53 */
            {8'h00}, /* 0x9f52 */
            {8'h00}, /* 0x9f51 */
            {8'h00}, /* 0x9f50 */
            {8'h00}, /* 0x9f4f */
            {8'h00}, /* 0x9f4e */
            {8'h00}, /* 0x9f4d */
            {8'h00}, /* 0x9f4c */
            {8'h00}, /* 0x9f4b */
            {8'h00}, /* 0x9f4a */
            {8'h00}, /* 0x9f49 */
            {8'h00}, /* 0x9f48 */
            {8'h00}, /* 0x9f47 */
            {8'h00}, /* 0x9f46 */
            {8'h00}, /* 0x9f45 */
            {8'h00}, /* 0x9f44 */
            {8'h00}, /* 0x9f43 */
            {8'h00}, /* 0x9f42 */
            {8'h00}, /* 0x9f41 */
            {8'h00}, /* 0x9f40 */
            {8'h00}, /* 0x9f3f */
            {8'h00}, /* 0x9f3e */
            {8'h00}, /* 0x9f3d */
            {8'h00}, /* 0x9f3c */
            {8'h00}, /* 0x9f3b */
            {8'h00}, /* 0x9f3a */
            {8'h00}, /* 0x9f39 */
            {8'h00}, /* 0x9f38 */
            {8'h00}, /* 0x9f37 */
            {8'h00}, /* 0x9f36 */
            {8'h00}, /* 0x9f35 */
            {8'h00}, /* 0x9f34 */
            {8'h00}, /* 0x9f33 */
            {8'h00}, /* 0x9f32 */
            {8'h00}, /* 0x9f31 */
            {8'h00}, /* 0x9f30 */
            {8'h00}, /* 0x9f2f */
            {8'h00}, /* 0x9f2e */
            {8'h00}, /* 0x9f2d */
            {8'h00}, /* 0x9f2c */
            {8'h00}, /* 0x9f2b */
            {8'h00}, /* 0x9f2a */
            {8'h00}, /* 0x9f29 */
            {8'h00}, /* 0x9f28 */
            {8'h00}, /* 0x9f27 */
            {8'h00}, /* 0x9f26 */
            {8'h00}, /* 0x9f25 */
            {8'h00}, /* 0x9f24 */
            {8'h00}, /* 0x9f23 */
            {8'h00}, /* 0x9f22 */
            {8'h00}, /* 0x9f21 */
            {8'h00}, /* 0x9f20 */
            {8'h00}, /* 0x9f1f */
            {8'h00}, /* 0x9f1e */
            {8'h00}, /* 0x9f1d */
            {8'h00}, /* 0x9f1c */
            {8'h00}, /* 0x9f1b */
            {8'h00}, /* 0x9f1a */
            {8'h00}, /* 0x9f19 */
            {8'h00}, /* 0x9f18 */
            {8'h00}, /* 0x9f17 */
            {8'h00}, /* 0x9f16 */
            {8'h00}, /* 0x9f15 */
            {8'h00}, /* 0x9f14 */
            {8'h00}, /* 0x9f13 */
            {8'h00}, /* 0x9f12 */
            {8'h00}, /* 0x9f11 */
            {8'h00}, /* 0x9f10 */
            {8'h00}, /* 0x9f0f */
            {8'h00}, /* 0x9f0e */
            {8'h00}, /* 0x9f0d */
            {8'h00}, /* 0x9f0c */
            {8'h00}, /* 0x9f0b */
            {8'h00}, /* 0x9f0a */
            {8'h00}, /* 0x9f09 */
            {8'h00}, /* 0x9f08 */
            {8'h00}, /* 0x9f07 */
            {8'h00}, /* 0x9f06 */
            {8'h00}, /* 0x9f05 */
            {8'h00}, /* 0x9f04 */
            {8'h00}, /* 0x9f03 */
            {8'h00}, /* 0x9f02 */
            {8'h00}, /* 0x9f01 */
            {8'h00}, /* 0x9f00 */
            {8'h00}, /* 0x9eff */
            {8'h00}, /* 0x9efe */
            {8'h00}, /* 0x9efd */
            {8'h00}, /* 0x9efc */
            {8'h00}, /* 0x9efb */
            {8'h00}, /* 0x9efa */
            {8'h00}, /* 0x9ef9 */
            {8'h00}, /* 0x9ef8 */
            {8'h00}, /* 0x9ef7 */
            {8'h00}, /* 0x9ef6 */
            {8'h00}, /* 0x9ef5 */
            {8'h00}, /* 0x9ef4 */
            {8'h00}, /* 0x9ef3 */
            {8'h00}, /* 0x9ef2 */
            {8'h00}, /* 0x9ef1 */
            {8'h00}, /* 0x9ef0 */
            {8'h00}, /* 0x9eef */
            {8'h00}, /* 0x9eee */
            {8'h00}, /* 0x9eed */
            {8'h00}, /* 0x9eec */
            {8'h00}, /* 0x9eeb */
            {8'h00}, /* 0x9eea */
            {8'h00}, /* 0x9ee9 */
            {8'h00}, /* 0x9ee8 */
            {8'h00}, /* 0x9ee7 */
            {8'h00}, /* 0x9ee6 */
            {8'h00}, /* 0x9ee5 */
            {8'h00}, /* 0x9ee4 */
            {8'h00}, /* 0x9ee3 */
            {8'h00}, /* 0x9ee2 */
            {8'h00}, /* 0x9ee1 */
            {8'h00}, /* 0x9ee0 */
            {8'h00}, /* 0x9edf */
            {8'h00}, /* 0x9ede */
            {8'h00}, /* 0x9edd */
            {8'h00}, /* 0x9edc */
            {8'h00}, /* 0x9edb */
            {8'h00}, /* 0x9eda */
            {8'h00}, /* 0x9ed9 */
            {8'h00}, /* 0x9ed8 */
            {8'h00}, /* 0x9ed7 */
            {8'h00}, /* 0x9ed6 */
            {8'h00}, /* 0x9ed5 */
            {8'h00}, /* 0x9ed4 */
            {8'h00}, /* 0x9ed3 */
            {8'h00}, /* 0x9ed2 */
            {8'h00}, /* 0x9ed1 */
            {8'h00}, /* 0x9ed0 */
            {8'h00}, /* 0x9ecf */
            {8'h00}, /* 0x9ece */
            {8'h00}, /* 0x9ecd */
            {8'h00}, /* 0x9ecc */
            {8'h00}, /* 0x9ecb */
            {8'h00}, /* 0x9eca */
            {8'h00}, /* 0x9ec9 */
            {8'h00}, /* 0x9ec8 */
            {8'h00}, /* 0x9ec7 */
            {8'h00}, /* 0x9ec6 */
            {8'h00}, /* 0x9ec5 */
            {8'h00}, /* 0x9ec4 */
            {8'h00}, /* 0x9ec3 */
            {8'h00}, /* 0x9ec2 */
            {8'h00}, /* 0x9ec1 */
            {8'h00}, /* 0x9ec0 */
            {8'h00}, /* 0x9ebf */
            {8'h00}, /* 0x9ebe */
            {8'h00}, /* 0x9ebd */
            {8'h00}, /* 0x9ebc */
            {8'h00}, /* 0x9ebb */
            {8'h00}, /* 0x9eba */
            {8'h00}, /* 0x9eb9 */
            {8'h00}, /* 0x9eb8 */
            {8'h00}, /* 0x9eb7 */
            {8'h00}, /* 0x9eb6 */
            {8'h00}, /* 0x9eb5 */
            {8'h00}, /* 0x9eb4 */
            {8'h00}, /* 0x9eb3 */
            {8'h00}, /* 0x9eb2 */
            {8'h00}, /* 0x9eb1 */
            {8'h00}, /* 0x9eb0 */
            {8'h00}, /* 0x9eaf */
            {8'h00}, /* 0x9eae */
            {8'h00}, /* 0x9ead */
            {8'h00}, /* 0x9eac */
            {8'h00}, /* 0x9eab */
            {8'h00}, /* 0x9eaa */
            {8'h00}, /* 0x9ea9 */
            {8'h00}, /* 0x9ea8 */
            {8'h00}, /* 0x9ea7 */
            {8'h00}, /* 0x9ea6 */
            {8'h00}, /* 0x9ea5 */
            {8'h00}, /* 0x9ea4 */
            {8'h00}, /* 0x9ea3 */
            {8'h00}, /* 0x9ea2 */
            {8'h00}, /* 0x9ea1 */
            {8'h00}, /* 0x9ea0 */
            {8'h00}, /* 0x9e9f */
            {8'h00}, /* 0x9e9e */
            {8'h00}, /* 0x9e9d */
            {8'h00}, /* 0x9e9c */
            {8'h00}, /* 0x9e9b */
            {8'h00}, /* 0x9e9a */
            {8'h00}, /* 0x9e99 */
            {8'h00}, /* 0x9e98 */
            {8'h00}, /* 0x9e97 */
            {8'h00}, /* 0x9e96 */
            {8'h00}, /* 0x9e95 */
            {8'h00}, /* 0x9e94 */
            {8'h00}, /* 0x9e93 */
            {8'h00}, /* 0x9e92 */
            {8'h00}, /* 0x9e91 */
            {8'h00}, /* 0x9e90 */
            {8'h00}, /* 0x9e8f */
            {8'h00}, /* 0x9e8e */
            {8'h00}, /* 0x9e8d */
            {8'h00}, /* 0x9e8c */
            {8'h00}, /* 0x9e8b */
            {8'h00}, /* 0x9e8a */
            {8'h00}, /* 0x9e89 */
            {8'h00}, /* 0x9e88 */
            {8'h00}, /* 0x9e87 */
            {8'h00}, /* 0x9e86 */
            {8'h00}, /* 0x9e85 */
            {8'h00}, /* 0x9e84 */
            {8'h00}, /* 0x9e83 */
            {8'h00}, /* 0x9e82 */
            {8'h00}, /* 0x9e81 */
            {8'h00}, /* 0x9e80 */
            {8'h00}, /* 0x9e7f */
            {8'h00}, /* 0x9e7e */
            {8'h00}, /* 0x9e7d */
            {8'h00}, /* 0x9e7c */
            {8'h00}, /* 0x9e7b */
            {8'h00}, /* 0x9e7a */
            {8'h00}, /* 0x9e79 */
            {8'h00}, /* 0x9e78 */
            {8'h00}, /* 0x9e77 */
            {8'h00}, /* 0x9e76 */
            {8'h00}, /* 0x9e75 */
            {8'h00}, /* 0x9e74 */
            {8'h00}, /* 0x9e73 */
            {8'h00}, /* 0x9e72 */
            {8'h00}, /* 0x9e71 */
            {8'h00}, /* 0x9e70 */
            {8'h00}, /* 0x9e6f */
            {8'h00}, /* 0x9e6e */
            {8'h00}, /* 0x9e6d */
            {8'h00}, /* 0x9e6c */
            {8'h00}, /* 0x9e6b */
            {8'h00}, /* 0x9e6a */
            {8'h00}, /* 0x9e69 */
            {8'h00}, /* 0x9e68 */
            {8'h00}, /* 0x9e67 */
            {8'h00}, /* 0x9e66 */
            {8'h00}, /* 0x9e65 */
            {8'h00}, /* 0x9e64 */
            {8'h00}, /* 0x9e63 */
            {8'h00}, /* 0x9e62 */
            {8'h00}, /* 0x9e61 */
            {8'h00}, /* 0x9e60 */
            {8'h00}, /* 0x9e5f */
            {8'h00}, /* 0x9e5e */
            {8'h00}, /* 0x9e5d */
            {8'h00}, /* 0x9e5c */
            {8'h00}, /* 0x9e5b */
            {8'h00}, /* 0x9e5a */
            {8'h00}, /* 0x9e59 */
            {8'h00}, /* 0x9e58 */
            {8'h00}, /* 0x9e57 */
            {8'h00}, /* 0x9e56 */
            {8'h00}, /* 0x9e55 */
            {8'h00}, /* 0x9e54 */
            {8'h00}, /* 0x9e53 */
            {8'h00}, /* 0x9e52 */
            {8'h00}, /* 0x9e51 */
            {8'h00}, /* 0x9e50 */
            {8'h00}, /* 0x9e4f */
            {8'h00}, /* 0x9e4e */
            {8'h00}, /* 0x9e4d */
            {8'h00}, /* 0x9e4c */
            {8'h00}, /* 0x9e4b */
            {8'h00}, /* 0x9e4a */
            {8'h00}, /* 0x9e49 */
            {8'h00}, /* 0x9e48 */
            {8'h00}, /* 0x9e47 */
            {8'h00}, /* 0x9e46 */
            {8'h00}, /* 0x9e45 */
            {8'h00}, /* 0x9e44 */
            {8'h00}, /* 0x9e43 */
            {8'h00}, /* 0x9e42 */
            {8'h00}, /* 0x9e41 */
            {8'h00}, /* 0x9e40 */
            {8'h00}, /* 0x9e3f */
            {8'h00}, /* 0x9e3e */
            {8'h00}, /* 0x9e3d */
            {8'h00}, /* 0x9e3c */
            {8'h00}, /* 0x9e3b */
            {8'h00}, /* 0x9e3a */
            {8'h00}, /* 0x9e39 */
            {8'h00}, /* 0x9e38 */
            {8'h00}, /* 0x9e37 */
            {8'h00}, /* 0x9e36 */
            {8'h00}, /* 0x9e35 */
            {8'h00}, /* 0x9e34 */
            {8'h00}, /* 0x9e33 */
            {8'h00}, /* 0x9e32 */
            {8'h00}, /* 0x9e31 */
            {8'h00}, /* 0x9e30 */
            {8'h00}, /* 0x9e2f */
            {8'h00}, /* 0x9e2e */
            {8'h00}, /* 0x9e2d */
            {8'h00}, /* 0x9e2c */
            {8'h00}, /* 0x9e2b */
            {8'h00}, /* 0x9e2a */
            {8'h00}, /* 0x9e29 */
            {8'h00}, /* 0x9e28 */
            {8'h00}, /* 0x9e27 */
            {8'h00}, /* 0x9e26 */
            {8'h00}, /* 0x9e25 */
            {8'h00}, /* 0x9e24 */
            {8'h00}, /* 0x9e23 */
            {8'h00}, /* 0x9e22 */
            {8'h00}, /* 0x9e21 */
            {8'h00}, /* 0x9e20 */
            {8'h00}, /* 0x9e1f */
            {8'h00}, /* 0x9e1e */
            {8'h00}, /* 0x9e1d */
            {8'h00}, /* 0x9e1c */
            {8'h00}, /* 0x9e1b */
            {8'h00}, /* 0x9e1a */
            {8'h00}, /* 0x9e19 */
            {8'h00}, /* 0x9e18 */
            {8'h00}, /* 0x9e17 */
            {8'h00}, /* 0x9e16 */
            {8'h00}, /* 0x9e15 */
            {8'h00}, /* 0x9e14 */
            {8'h00}, /* 0x9e13 */
            {8'h00}, /* 0x9e12 */
            {8'h00}, /* 0x9e11 */
            {8'h00}, /* 0x9e10 */
            {8'h00}, /* 0x9e0f */
            {8'h00}, /* 0x9e0e */
            {8'h00}, /* 0x9e0d */
            {8'h00}, /* 0x9e0c */
            {8'h00}, /* 0x9e0b */
            {8'h00}, /* 0x9e0a */
            {8'h00}, /* 0x9e09 */
            {8'h00}, /* 0x9e08 */
            {8'h00}, /* 0x9e07 */
            {8'h00}, /* 0x9e06 */
            {8'h00}, /* 0x9e05 */
            {8'h00}, /* 0x9e04 */
            {8'h00}, /* 0x9e03 */
            {8'h00}, /* 0x9e02 */
            {8'h00}, /* 0x9e01 */
            {8'h00}, /* 0x9e00 */
            {8'h00}, /* 0x9dff */
            {8'h00}, /* 0x9dfe */
            {8'h00}, /* 0x9dfd */
            {8'h00}, /* 0x9dfc */
            {8'h00}, /* 0x9dfb */
            {8'h00}, /* 0x9dfa */
            {8'h00}, /* 0x9df9 */
            {8'h00}, /* 0x9df8 */
            {8'h00}, /* 0x9df7 */
            {8'h00}, /* 0x9df6 */
            {8'h00}, /* 0x9df5 */
            {8'h00}, /* 0x9df4 */
            {8'h00}, /* 0x9df3 */
            {8'h00}, /* 0x9df2 */
            {8'h00}, /* 0x9df1 */
            {8'h00}, /* 0x9df0 */
            {8'h00}, /* 0x9def */
            {8'h00}, /* 0x9dee */
            {8'h00}, /* 0x9ded */
            {8'h00}, /* 0x9dec */
            {8'h00}, /* 0x9deb */
            {8'h00}, /* 0x9dea */
            {8'h00}, /* 0x9de9 */
            {8'h00}, /* 0x9de8 */
            {8'h00}, /* 0x9de7 */
            {8'h00}, /* 0x9de6 */
            {8'h00}, /* 0x9de5 */
            {8'h00}, /* 0x9de4 */
            {8'h00}, /* 0x9de3 */
            {8'h00}, /* 0x9de2 */
            {8'h00}, /* 0x9de1 */
            {8'h00}, /* 0x9de0 */
            {8'h00}, /* 0x9ddf */
            {8'h00}, /* 0x9dde */
            {8'h00}, /* 0x9ddd */
            {8'h00}, /* 0x9ddc */
            {8'h00}, /* 0x9ddb */
            {8'h00}, /* 0x9dda */
            {8'h00}, /* 0x9dd9 */
            {8'h00}, /* 0x9dd8 */
            {8'h00}, /* 0x9dd7 */
            {8'h00}, /* 0x9dd6 */
            {8'h00}, /* 0x9dd5 */
            {8'h00}, /* 0x9dd4 */
            {8'h00}, /* 0x9dd3 */
            {8'h00}, /* 0x9dd2 */
            {8'h00}, /* 0x9dd1 */
            {8'h00}, /* 0x9dd0 */
            {8'h00}, /* 0x9dcf */
            {8'h00}, /* 0x9dce */
            {8'h00}, /* 0x9dcd */
            {8'h00}, /* 0x9dcc */
            {8'h00}, /* 0x9dcb */
            {8'h00}, /* 0x9dca */
            {8'h00}, /* 0x9dc9 */
            {8'h00}, /* 0x9dc8 */
            {8'h00}, /* 0x9dc7 */
            {8'h00}, /* 0x9dc6 */
            {8'h00}, /* 0x9dc5 */
            {8'h00}, /* 0x9dc4 */
            {8'h00}, /* 0x9dc3 */
            {8'h00}, /* 0x9dc2 */
            {8'h00}, /* 0x9dc1 */
            {8'h00}, /* 0x9dc0 */
            {8'h00}, /* 0x9dbf */
            {8'h00}, /* 0x9dbe */
            {8'h00}, /* 0x9dbd */
            {8'h00}, /* 0x9dbc */
            {8'h00}, /* 0x9dbb */
            {8'h00}, /* 0x9dba */
            {8'h00}, /* 0x9db9 */
            {8'h00}, /* 0x9db8 */
            {8'h00}, /* 0x9db7 */
            {8'h00}, /* 0x9db6 */
            {8'h00}, /* 0x9db5 */
            {8'h00}, /* 0x9db4 */
            {8'h00}, /* 0x9db3 */
            {8'h00}, /* 0x9db2 */
            {8'h00}, /* 0x9db1 */
            {8'h00}, /* 0x9db0 */
            {8'h00}, /* 0x9daf */
            {8'h00}, /* 0x9dae */
            {8'h00}, /* 0x9dad */
            {8'h00}, /* 0x9dac */
            {8'h00}, /* 0x9dab */
            {8'h00}, /* 0x9daa */
            {8'h00}, /* 0x9da9 */
            {8'h00}, /* 0x9da8 */
            {8'h00}, /* 0x9da7 */
            {8'h00}, /* 0x9da6 */
            {8'h00}, /* 0x9da5 */
            {8'h00}, /* 0x9da4 */
            {8'h00}, /* 0x9da3 */
            {8'h00}, /* 0x9da2 */
            {8'h00}, /* 0x9da1 */
            {8'h00}, /* 0x9da0 */
            {8'h00}, /* 0x9d9f */
            {8'h00}, /* 0x9d9e */
            {8'h00}, /* 0x9d9d */
            {8'h00}, /* 0x9d9c */
            {8'h00}, /* 0x9d9b */
            {8'h00}, /* 0x9d9a */
            {8'h00}, /* 0x9d99 */
            {8'h00}, /* 0x9d98 */
            {8'h00}, /* 0x9d97 */
            {8'h00}, /* 0x9d96 */
            {8'h00}, /* 0x9d95 */
            {8'h00}, /* 0x9d94 */
            {8'h00}, /* 0x9d93 */
            {8'h00}, /* 0x9d92 */
            {8'h00}, /* 0x9d91 */
            {8'h00}, /* 0x9d90 */
            {8'h00}, /* 0x9d8f */
            {8'h00}, /* 0x9d8e */
            {8'h00}, /* 0x9d8d */
            {8'h00}, /* 0x9d8c */
            {8'h00}, /* 0x9d8b */
            {8'h00}, /* 0x9d8a */
            {8'h00}, /* 0x9d89 */
            {8'h00}, /* 0x9d88 */
            {8'h00}, /* 0x9d87 */
            {8'h00}, /* 0x9d86 */
            {8'h00}, /* 0x9d85 */
            {8'h00}, /* 0x9d84 */
            {8'h00}, /* 0x9d83 */
            {8'h00}, /* 0x9d82 */
            {8'h00}, /* 0x9d81 */
            {8'h00}, /* 0x9d80 */
            {8'h00}, /* 0x9d7f */
            {8'h00}, /* 0x9d7e */
            {8'h00}, /* 0x9d7d */
            {8'h00}, /* 0x9d7c */
            {8'h00}, /* 0x9d7b */
            {8'h00}, /* 0x9d7a */
            {8'h00}, /* 0x9d79 */
            {8'h00}, /* 0x9d78 */
            {8'h00}, /* 0x9d77 */
            {8'h00}, /* 0x9d76 */
            {8'h00}, /* 0x9d75 */
            {8'h00}, /* 0x9d74 */
            {8'h00}, /* 0x9d73 */
            {8'h00}, /* 0x9d72 */
            {8'h00}, /* 0x9d71 */
            {8'h00}, /* 0x9d70 */
            {8'h00}, /* 0x9d6f */
            {8'h00}, /* 0x9d6e */
            {8'h00}, /* 0x9d6d */
            {8'h00}, /* 0x9d6c */
            {8'h00}, /* 0x9d6b */
            {8'h00}, /* 0x9d6a */
            {8'h00}, /* 0x9d69 */
            {8'h00}, /* 0x9d68 */
            {8'h00}, /* 0x9d67 */
            {8'h00}, /* 0x9d66 */
            {8'h00}, /* 0x9d65 */
            {8'h00}, /* 0x9d64 */
            {8'h00}, /* 0x9d63 */
            {8'h00}, /* 0x9d62 */
            {8'h00}, /* 0x9d61 */
            {8'h00}, /* 0x9d60 */
            {8'h00}, /* 0x9d5f */
            {8'h00}, /* 0x9d5e */
            {8'h00}, /* 0x9d5d */
            {8'h00}, /* 0x9d5c */
            {8'h00}, /* 0x9d5b */
            {8'h00}, /* 0x9d5a */
            {8'h00}, /* 0x9d59 */
            {8'h00}, /* 0x9d58 */
            {8'h00}, /* 0x9d57 */
            {8'h00}, /* 0x9d56 */
            {8'h00}, /* 0x9d55 */
            {8'h00}, /* 0x9d54 */
            {8'h00}, /* 0x9d53 */
            {8'h00}, /* 0x9d52 */
            {8'h00}, /* 0x9d51 */
            {8'h00}, /* 0x9d50 */
            {8'h00}, /* 0x9d4f */
            {8'h00}, /* 0x9d4e */
            {8'h00}, /* 0x9d4d */
            {8'h00}, /* 0x9d4c */
            {8'h00}, /* 0x9d4b */
            {8'h00}, /* 0x9d4a */
            {8'h00}, /* 0x9d49 */
            {8'h00}, /* 0x9d48 */
            {8'h00}, /* 0x9d47 */
            {8'h00}, /* 0x9d46 */
            {8'h00}, /* 0x9d45 */
            {8'h00}, /* 0x9d44 */
            {8'h00}, /* 0x9d43 */
            {8'h00}, /* 0x9d42 */
            {8'h00}, /* 0x9d41 */
            {8'h00}, /* 0x9d40 */
            {8'h00}, /* 0x9d3f */
            {8'h00}, /* 0x9d3e */
            {8'h00}, /* 0x9d3d */
            {8'h00}, /* 0x9d3c */
            {8'h00}, /* 0x9d3b */
            {8'h00}, /* 0x9d3a */
            {8'h00}, /* 0x9d39 */
            {8'h00}, /* 0x9d38 */
            {8'h00}, /* 0x9d37 */
            {8'h00}, /* 0x9d36 */
            {8'h00}, /* 0x9d35 */
            {8'h00}, /* 0x9d34 */
            {8'h00}, /* 0x9d33 */
            {8'h00}, /* 0x9d32 */
            {8'h00}, /* 0x9d31 */
            {8'h00}, /* 0x9d30 */
            {8'h00}, /* 0x9d2f */
            {8'h00}, /* 0x9d2e */
            {8'h00}, /* 0x9d2d */
            {8'h00}, /* 0x9d2c */
            {8'h00}, /* 0x9d2b */
            {8'h00}, /* 0x9d2a */
            {8'h00}, /* 0x9d29 */
            {8'h00}, /* 0x9d28 */
            {8'h00}, /* 0x9d27 */
            {8'h00}, /* 0x9d26 */
            {8'h00}, /* 0x9d25 */
            {8'h00}, /* 0x9d24 */
            {8'h00}, /* 0x9d23 */
            {8'h00}, /* 0x9d22 */
            {8'h00}, /* 0x9d21 */
            {8'h00}, /* 0x9d20 */
            {8'h00}, /* 0x9d1f */
            {8'h00}, /* 0x9d1e */
            {8'h00}, /* 0x9d1d */
            {8'h00}, /* 0x9d1c */
            {8'h00}, /* 0x9d1b */
            {8'h00}, /* 0x9d1a */
            {8'h00}, /* 0x9d19 */
            {8'h00}, /* 0x9d18 */
            {8'h00}, /* 0x9d17 */
            {8'h00}, /* 0x9d16 */
            {8'h00}, /* 0x9d15 */
            {8'h00}, /* 0x9d14 */
            {8'h00}, /* 0x9d13 */
            {8'h00}, /* 0x9d12 */
            {8'h00}, /* 0x9d11 */
            {8'h00}, /* 0x9d10 */
            {8'h00}, /* 0x9d0f */
            {8'h00}, /* 0x9d0e */
            {8'h00}, /* 0x9d0d */
            {8'h00}, /* 0x9d0c */
            {8'h00}, /* 0x9d0b */
            {8'h00}, /* 0x9d0a */
            {8'h00}, /* 0x9d09 */
            {8'h00}, /* 0x9d08 */
            {8'h00}, /* 0x9d07 */
            {8'h00}, /* 0x9d06 */
            {8'h00}, /* 0x9d05 */
            {8'h00}, /* 0x9d04 */
            {8'h00}, /* 0x9d03 */
            {8'h00}, /* 0x9d02 */
            {8'h00}, /* 0x9d01 */
            {8'h00}, /* 0x9d00 */
            {8'h00}, /* 0x9cff */
            {8'h00}, /* 0x9cfe */
            {8'h00}, /* 0x9cfd */
            {8'h00}, /* 0x9cfc */
            {8'h00}, /* 0x9cfb */
            {8'h00}, /* 0x9cfa */
            {8'h00}, /* 0x9cf9 */
            {8'h00}, /* 0x9cf8 */
            {8'h00}, /* 0x9cf7 */
            {8'h00}, /* 0x9cf6 */
            {8'h00}, /* 0x9cf5 */
            {8'h00}, /* 0x9cf4 */
            {8'h00}, /* 0x9cf3 */
            {8'h00}, /* 0x9cf2 */
            {8'h00}, /* 0x9cf1 */
            {8'h00}, /* 0x9cf0 */
            {8'h00}, /* 0x9cef */
            {8'h00}, /* 0x9cee */
            {8'h00}, /* 0x9ced */
            {8'h00}, /* 0x9cec */
            {8'h00}, /* 0x9ceb */
            {8'h00}, /* 0x9cea */
            {8'h00}, /* 0x9ce9 */
            {8'h00}, /* 0x9ce8 */
            {8'h00}, /* 0x9ce7 */
            {8'h00}, /* 0x9ce6 */
            {8'h00}, /* 0x9ce5 */
            {8'h00}, /* 0x9ce4 */
            {8'h00}, /* 0x9ce3 */
            {8'h00}, /* 0x9ce2 */
            {8'h00}, /* 0x9ce1 */
            {8'h00}, /* 0x9ce0 */
            {8'h00}, /* 0x9cdf */
            {8'h00}, /* 0x9cde */
            {8'h00}, /* 0x9cdd */
            {8'h00}, /* 0x9cdc */
            {8'h00}, /* 0x9cdb */
            {8'h00}, /* 0x9cda */
            {8'h00}, /* 0x9cd9 */
            {8'h00}, /* 0x9cd8 */
            {8'h00}, /* 0x9cd7 */
            {8'h00}, /* 0x9cd6 */
            {8'h00}, /* 0x9cd5 */
            {8'h00}, /* 0x9cd4 */
            {8'h00}, /* 0x9cd3 */
            {8'h00}, /* 0x9cd2 */
            {8'h00}, /* 0x9cd1 */
            {8'h00}, /* 0x9cd0 */
            {8'h00}, /* 0x9ccf */
            {8'h00}, /* 0x9cce */
            {8'h00}, /* 0x9ccd */
            {8'h00}, /* 0x9ccc */
            {8'h00}, /* 0x9ccb */
            {8'h00}, /* 0x9cca */
            {8'h00}, /* 0x9cc9 */
            {8'h00}, /* 0x9cc8 */
            {8'h00}, /* 0x9cc7 */
            {8'h00}, /* 0x9cc6 */
            {8'h00}, /* 0x9cc5 */
            {8'h00}, /* 0x9cc4 */
            {8'h00}, /* 0x9cc3 */
            {8'h00}, /* 0x9cc2 */
            {8'h00}, /* 0x9cc1 */
            {8'h00}, /* 0x9cc0 */
            {8'h00}, /* 0x9cbf */
            {8'h00}, /* 0x9cbe */
            {8'h00}, /* 0x9cbd */
            {8'h00}, /* 0x9cbc */
            {8'h00}, /* 0x9cbb */
            {8'h00}, /* 0x9cba */
            {8'h00}, /* 0x9cb9 */
            {8'h00}, /* 0x9cb8 */
            {8'h00}, /* 0x9cb7 */
            {8'h00}, /* 0x9cb6 */
            {8'h00}, /* 0x9cb5 */
            {8'h00}, /* 0x9cb4 */
            {8'h00}, /* 0x9cb3 */
            {8'h00}, /* 0x9cb2 */
            {8'h00}, /* 0x9cb1 */
            {8'h00}, /* 0x9cb0 */
            {8'h00}, /* 0x9caf */
            {8'h00}, /* 0x9cae */
            {8'h00}, /* 0x9cad */
            {8'h00}, /* 0x9cac */
            {8'h00}, /* 0x9cab */
            {8'h00}, /* 0x9caa */
            {8'h00}, /* 0x9ca9 */
            {8'h00}, /* 0x9ca8 */
            {8'h00}, /* 0x9ca7 */
            {8'h00}, /* 0x9ca6 */
            {8'h00}, /* 0x9ca5 */
            {8'h00}, /* 0x9ca4 */
            {8'h00}, /* 0x9ca3 */
            {8'h00}, /* 0x9ca2 */
            {8'h00}, /* 0x9ca1 */
            {8'h00}, /* 0x9ca0 */
            {8'h00}, /* 0x9c9f */
            {8'h00}, /* 0x9c9e */
            {8'h00}, /* 0x9c9d */
            {8'h00}, /* 0x9c9c */
            {8'h00}, /* 0x9c9b */
            {8'h00}, /* 0x9c9a */
            {8'h00}, /* 0x9c99 */
            {8'h00}, /* 0x9c98 */
            {8'h00}, /* 0x9c97 */
            {8'h00}, /* 0x9c96 */
            {8'h00}, /* 0x9c95 */
            {8'h00}, /* 0x9c94 */
            {8'h00}, /* 0x9c93 */
            {8'h00}, /* 0x9c92 */
            {8'h00}, /* 0x9c91 */
            {8'h00}, /* 0x9c90 */
            {8'h00}, /* 0x9c8f */
            {8'h00}, /* 0x9c8e */
            {8'h00}, /* 0x9c8d */
            {8'h00}, /* 0x9c8c */
            {8'h00}, /* 0x9c8b */
            {8'h00}, /* 0x9c8a */
            {8'h00}, /* 0x9c89 */
            {8'h00}, /* 0x9c88 */
            {8'h00}, /* 0x9c87 */
            {8'h00}, /* 0x9c86 */
            {8'h00}, /* 0x9c85 */
            {8'h00}, /* 0x9c84 */
            {8'h00}, /* 0x9c83 */
            {8'h00}, /* 0x9c82 */
            {8'h00}, /* 0x9c81 */
            {8'h00}, /* 0x9c80 */
            {8'h00}, /* 0x9c7f */
            {8'h00}, /* 0x9c7e */
            {8'h00}, /* 0x9c7d */
            {8'h00}, /* 0x9c7c */
            {8'h00}, /* 0x9c7b */
            {8'h00}, /* 0x9c7a */
            {8'h00}, /* 0x9c79 */
            {8'h00}, /* 0x9c78 */
            {8'h00}, /* 0x9c77 */
            {8'h00}, /* 0x9c76 */
            {8'h00}, /* 0x9c75 */
            {8'h00}, /* 0x9c74 */
            {8'h00}, /* 0x9c73 */
            {8'h00}, /* 0x9c72 */
            {8'h00}, /* 0x9c71 */
            {8'h00}, /* 0x9c70 */
            {8'h00}, /* 0x9c6f */
            {8'h00}, /* 0x9c6e */
            {8'h00}, /* 0x9c6d */
            {8'h00}, /* 0x9c6c */
            {8'h00}, /* 0x9c6b */
            {8'h00}, /* 0x9c6a */
            {8'h00}, /* 0x9c69 */
            {8'h00}, /* 0x9c68 */
            {8'h00}, /* 0x9c67 */
            {8'h00}, /* 0x9c66 */
            {8'h00}, /* 0x9c65 */
            {8'h00}, /* 0x9c64 */
            {8'h00}, /* 0x9c63 */
            {8'h00}, /* 0x9c62 */
            {8'h00}, /* 0x9c61 */
            {8'h00}, /* 0x9c60 */
            {8'h00}, /* 0x9c5f */
            {8'h00}, /* 0x9c5e */
            {8'h00}, /* 0x9c5d */
            {8'h00}, /* 0x9c5c */
            {8'h00}, /* 0x9c5b */
            {8'h00}, /* 0x9c5a */
            {8'h00}, /* 0x9c59 */
            {8'h00}, /* 0x9c58 */
            {8'h00}, /* 0x9c57 */
            {8'h00}, /* 0x9c56 */
            {8'h00}, /* 0x9c55 */
            {8'h00}, /* 0x9c54 */
            {8'h00}, /* 0x9c53 */
            {8'h00}, /* 0x9c52 */
            {8'h00}, /* 0x9c51 */
            {8'h00}, /* 0x9c50 */
            {8'h00}, /* 0x9c4f */
            {8'h00}, /* 0x9c4e */
            {8'h00}, /* 0x9c4d */
            {8'h00}, /* 0x9c4c */
            {8'h00}, /* 0x9c4b */
            {8'h00}, /* 0x9c4a */
            {8'h00}, /* 0x9c49 */
            {8'h00}, /* 0x9c48 */
            {8'h00}, /* 0x9c47 */
            {8'h00}, /* 0x9c46 */
            {8'h00}, /* 0x9c45 */
            {8'h00}, /* 0x9c44 */
            {8'h00}, /* 0x9c43 */
            {8'h00}, /* 0x9c42 */
            {8'h00}, /* 0x9c41 */
            {8'h00}, /* 0x9c40 */
            {8'h00}, /* 0x9c3f */
            {8'h00}, /* 0x9c3e */
            {8'h00}, /* 0x9c3d */
            {8'h00}, /* 0x9c3c */
            {8'h00}, /* 0x9c3b */
            {8'h00}, /* 0x9c3a */
            {8'h00}, /* 0x9c39 */
            {8'h00}, /* 0x9c38 */
            {8'h00}, /* 0x9c37 */
            {8'h00}, /* 0x9c36 */
            {8'h00}, /* 0x9c35 */
            {8'h00}, /* 0x9c34 */
            {8'h00}, /* 0x9c33 */
            {8'h00}, /* 0x9c32 */
            {8'h00}, /* 0x9c31 */
            {8'h00}, /* 0x9c30 */
            {8'h00}, /* 0x9c2f */
            {8'h00}, /* 0x9c2e */
            {8'h00}, /* 0x9c2d */
            {8'h00}, /* 0x9c2c */
            {8'h00}, /* 0x9c2b */
            {8'h00}, /* 0x9c2a */
            {8'h00}, /* 0x9c29 */
            {8'h00}, /* 0x9c28 */
            {8'h00}, /* 0x9c27 */
            {8'h00}, /* 0x9c26 */
            {8'h00}, /* 0x9c25 */
            {8'h00}, /* 0x9c24 */
            {8'h00}, /* 0x9c23 */
            {8'h00}, /* 0x9c22 */
            {8'h00}, /* 0x9c21 */
            {8'h00}, /* 0x9c20 */
            {8'h00}, /* 0x9c1f */
            {8'h00}, /* 0x9c1e */
            {8'h00}, /* 0x9c1d */
            {8'h00}, /* 0x9c1c */
            {8'h00}, /* 0x9c1b */
            {8'h00}, /* 0x9c1a */
            {8'h00}, /* 0x9c19 */
            {8'h00}, /* 0x9c18 */
            {8'h00}, /* 0x9c17 */
            {8'h00}, /* 0x9c16 */
            {8'h00}, /* 0x9c15 */
            {8'h00}, /* 0x9c14 */
            {8'h00}, /* 0x9c13 */
            {8'h00}, /* 0x9c12 */
            {8'h00}, /* 0x9c11 */
            {8'h00}, /* 0x9c10 */
            {8'h00}, /* 0x9c0f */
            {8'h00}, /* 0x9c0e */
            {8'h00}, /* 0x9c0d */
            {8'h00}, /* 0x9c0c */
            {8'h00}, /* 0x9c0b */
            {8'h00}, /* 0x9c0a */
            {8'h00}, /* 0x9c09 */
            {8'h00}, /* 0x9c08 */
            {8'h00}, /* 0x9c07 */
            {8'h00}, /* 0x9c06 */
            {8'h00}, /* 0x9c05 */
            {8'h00}, /* 0x9c04 */
            {8'h00}, /* 0x9c03 */
            {8'h00}, /* 0x9c02 */
            {8'h00}, /* 0x9c01 */
            {8'h00}, /* 0x9c00 */
            {8'h00}, /* 0x9bff */
            {8'h00}, /* 0x9bfe */
            {8'h00}, /* 0x9bfd */
            {8'h00}, /* 0x9bfc */
            {8'h00}, /* 0x9bfb */
            {8'h00}, /* 0x9bfa */
            {8'h00}, /* 0x9bf9 */
            {8'h00}, /* 0x9bf8 */
            {8'h00}, /* 0x9bf7 */
            {8'h00}, /* 0x9bf6 */
            {8'h00}, /* 0x9bf5 */
            {8'h00}, /* 0x9bf4 */
            {8'h00}, /* 0x9bf3 */
            {8'h00}, /* 0x9bf2 */
            {8'h00}, /* 0x9bf1 */
            {8'h00}, /* 0x9bf0 */
            {8'h00}, /* 0x9bef */
            {8'h00}, /* 0x9bee */
            {8'h00}, /* 0x9bed */
            {8'h00}, /* 0x9bec */
            {8'h00}, /* 0x9beb */
            {8'h00}, /* 0x9bea */
            {8'h00}, /* 0x9be9 */
            {8'h00}, /* 0x9be8 */
            {8'h00}, /* 0x9be7 */
            {8'h00}, /* 0x9be6 */
            {8'h00}, /* 0x9be5 */
            {8'h00}, /* 0x9be4 */
            {8'h00}, /* 0x9be3 */
            {8'h00}, /* 0x9be2 */
            {8'h00}, /* 0x9be1 */
            {8'h00}, /* 0x9be0 */
            {8'h00}, /* 0x9bdf */
            {8'h00}, /* 0x9bde */
            {8'h00}, /* 0x9bdd */
            {8'h00}, /* 0x9bdc */
            {8'h00}, /* 0x9bdb */
            {8'h00}, /* 0x9bda */
            {8'h00}, /* 0x9bd9 */
            {8'h00}, /* 0x9bd8 */
            {8'h00}, /* 0x9bd7 */
            {8'h00}, /* 0x9bd6 */
            {8'h00}, /* 0x9bd5 */
            {8'h00}, /* 0x9bd4 */
            {8'h00}, /* 0x9bd3 */
            {8'h00}, /* 0x9bd2 */
            {8'h00}, /* 0x9bd1 */
            {8'h00}, /* 0x9bd0 */
            {8'h00}, /* 0x9bcf */
            {8'h00}, /* 0x9bce */
            {8'h00}, /* 0x9bcd */
            {8'h00}, /* 0x9bcc */
            {8'h00}, /* 0x9bcb */
            {8'h00}, /* 0x9bca */
            {8'h00}, /* 0x9bc9 */
            {8'h00}, /* 0x9bc8 */
            {8'h00}, /* 0x9bc7 */
            {8'h00}, /* 0x9bc6 */
            {8'h00}, /* 0x9bc5 */
            {8'h00}, /* 0x9bc4 */
            {8'h00}, /* 0x9bc3 */
            {8'h00}, /* 0x9bc2 */
            {8'h00}, /* 0x9bc1 */
            {8'h00}, /* 0x9bc0 */
            {8'h00}, /* 0x9bbf */
            {8'h00}, /* 0x9bbe */
            {8'h00}, /* 0x9bbd */
            {8'h00}, /* 0x9bbc */
            {8'h00}, /* 0x9bbb */
            {8'h00}, /* 0x9bba */
            {8'h00}, /* 0x9bb9 */
            {8'h00}, /* 0x9bb8 */
            {8'h00}, /* 0x9bb7 */
            {8'h00}, /* 0x9bb6 */
            {8'h00}, /* 0x9bb5 */
            {8'h00}, /* 0x9bb4 */
            {8'h00}, /* 0x9bb3 */
            {8'h00}, /* 0x9bb2 */
            {8'h00}, /* 0x9bb1 */
            {8'h00}, /* 0x9bb0 */
            {8'h00}, /* 0x9baf */
            {8'h00}, /* 0x9bae */
            {8'h00}, /* 0x9bad */
            {8'h00}, /* 0x9bac */
            {8'h00}, /* 0x9bab */
            {8'h00}, /* 0x9baa */
            {8'h00}, /* 0x9ba9 */
            {8'h00}, /* 0x9ba8 */
            {8'h00}, /* 0x9ba7 */
            {8'h00}, /* 0x9ba6 */
            {8'h00}, /* 0x9ba5 */
            {8'h00}, /* 0x9ba4 */
            {8'h00}, /* 0x9ba3 */
            {8'h00}, /* 0x9ba2 */
            {8'h00}, /* 0x9ba1 */
            {8'h00}, /* 0x9ba0 */
            {8'h00}, /* 0x9b9f */
            {8'h00}, /* 0x9b9e */
            {8'h00}, /* 0x9b9d */
            {8'h00}, /* 0x9b9c */
            {8'h00}, /* 0x9b9b */
            {8'h00}, /* 0x9b9a */
            {8'h00}, /* 0x9b99 */
            {8'h00}, /* 0x9b98 */
            {8'h00}, /* 0x9b97 */
            {8'h00}, /* 0x9b96 */
            {8'h00}, /* 0x9b95 */
            {8'h00}, /* 0x9b94 */
            {8'h00}, /* 0x9b93 */
            {8'h00}, /* 0x9b92 */
            {8'h00}, /* 0x9b91 */
            {8'h00}, /* 0x9b90 */
            {8'h00}, /* 0x9b8f */
            {8'h00}, /* 0x9b8e */
            {8'h00}, /* 0x9b8d */
            {8'h00}, /* 0x9b8c */
            {8'h00}, /* 0x9b8b */
            {8'h00}, /* 0x9b8a */
            {8'h00}, /* 0x9b89 */
            {8'h00}, /* 0x9b88 */
            {8'h00}, /* 0x9b87 */
            {8'h00}, /* 0x9b86 */
            {8'h00}, /* 0x9b85 */
            {8'h00}, /* 0x9b84 */
            {8'h00}, /* 0x9b83 */
            {8'h00}, /* 0x9b82 */
            {8'h00}, /* 0x9b81 */
            {8'h00}, /* 0x9b80 */
            {8'h00}, /* 0x9b7f */
            {8'h00}, /* 0x9b7e */
            {8'h00}, /* 0x9b7d */
            {8'h00}, /* 0x9b7c */
            {8'h00}, /* 0x9b7b */
            {8'h00}, /* 0x9b7a */
            {8'h00}, /* 0x9b79 */
            {8'h00}, /* 0x9b78 */
            {8'h00}, /* 0x9b77 */
            {8'h00}, /* 0x9b76 */
            {8'h00}, /* 0x9b75 */
            {8'h00}, /* 0x9b74 */
            {8'h00}, /* 0x9b73 */
            {8'h00}, /* 0x9b72 */
            {8'h00}, /* 0x9b71 */
            {8'h00}, /* 0x9b70 */
            {8'h00}, /* 0x9b6f */
            {8'h00}, /* 0x9b6e */
            {8'h00}, /* 0x9b6d */
            {8'h00}, /* 0x9b6c */
            {8'h00}, /* 0x9b6b */
            {8'h00}, /* 0x9b6a */
            {8'h00}, /* 0x9b69 */
            {8'h00}, /* 0x9b68 */
            {8'h00}, /* 0x9b67 */
            {8'h00}, /* 0x9b66 */
            {8'h00}, /* 0x9b65 */
            {8'h00}, /* 0x9b64 */
            {8'h00}, /* 0x9b63 */
            {8'h00}, /* 0x9b62 */
            {8'h00}, /* 0x9b61 */
            {8'h00}, /* 0x9b60 */
            {8'h00}, /* 0x9b5f */
            {8'h00}, /* 0x9b5e */
            {8'h00}, /* 0x9b5d */
            {8'h00}, /* 0x9b5c */
            {8'h00}, /* 0x9b5b */
            {8'h00}, /* 0x9b5a */
            {8'h00}, /* 0x9b59 */
            {8'h00}, /* 0x9b58 */
            {8'h00}, /* 0x9b57 */
            {8'h00}, /* 0x9b56 */
            {8'h00}, /* 0x9b55 */
            {8'h00}, /* 0x9b54 */
            {8'h00}, /* 0x9b53 */
            {8'h00}, /* 0x9b52 */
            {8'h00}, /* 0x9b51 */
            {8'h00}, /* 0x9b50 */
            {8'h00}, /* 0x9b4f */
            {8'h00}, /* 0x9b4e */
            {8'h00}, /* 0x9b4d */
            {8'h00}, /* 0x9b4c */
            {8'h00}, /* 0x9b4b */
            {8'h00}, /* 0x9b4a */
            {8'h00}, /* 0x9b49 */
            {8'h00}, /* 0x9b48 */
            {8'h00}, /* 0x9b47 */
            {8'h00}, /* 0x9b46 */
            {8'h00}, /* 0x9b45 */
            {8'h00}, /* 0x9b44 */
            {8'h00}, /* 0x9b43 */
            {8'h00}, /* 0x9b42 */
            {8'h00}, /* 0x9b41 */
            {8'h00}, /* 0x9b40 */
            {8'h00}, /* 0x9b3f */
            {8'h00}, /* 0x9b3e */
            {8'h00}, /* 0x9b3d */
            {8'h00}, /* 0x9b3c */
            {8'h00}, /* 0x9b3b */
            {8'h00}, /* 0x9b3a */
            {8'h00}, /* 0x9b39 */
            {8'h00}, /* 0x9b38 */
            {8'h00}, /* 0x9b37 */
            {8'h00}, /* 0x9b36 */
            {8'h00}, /* 0x9b35 */
            {8'h00}, /* 0x9b34 */
            {8'h00}, /* 0x9b33 */
            {8'h00}, /* 0x9b32 */
            {8'h00}, /* 0x9b31 */
            {8'h00}, /* 0x9b30 */
            {8'h00}, /* 0x9b2f */
            {8'h00}, /* 0x9b2e */
            {8'h00}, /* 0x9b2d */
            {8'h00}, /* 0x9b2c */
            {8'h00}, /* 0x9b2b */
            {8'h00}, /* 0x9b2a */
            {8'h00}, /* 0x9b29 */
            {8'h00}, /* 0x9b28 */
            {8'h00}, /* 0x9b27 */
            {8'h00}, /* 0x9b26 */
            {8'h00}, /* 0x9b25 */
            {8'h00}, /* 0x9b24 */
            {8'h00}, /* 0x9b23 */
            {8'h00}, /* 0x9b22 */
            {8'h00}, /* 0x9b21 */
            {8'h00}, /* 0x9b20 */
            {8'h00}, /* 0x9b1f */
            {8'h00}, /* 0x9b1e */
            {8'h00}, /* 0x9b1d */
            {8'h00}, /* 0x9b1c */
            {8'h00}, /* 0x9b1b */
            {8'h00}, /* 0x9b1a */
            {8'h00}, /* 0x9b19 */
            {8'h00}, /* 0x9b18 */
            {8'h00}, /* 0x9b17 */
            {8'h00}, /* 0x9b16 */
            {8'h00}, /* 0x9b15 */
            {8'h00}, /* 0x9b14 */
            {8'h00}, /* 0x9b13 */
            {8'h00}, /* 0x9b12 */
            {8'h00}, /* 0x9b11 */
            {8'h00}, /* 0x9b10 */
            {8'h00}, /* 0x9b0f */
            {8'h00}, /* 0x9b0e */
            {8'h00}, /* 0x9b0d */
            {8'h00}, /* 0x9b0c */
            {8'h00}, /* 0x9b0b */
            {8'h00}, /* 0x9b0a */
            {8'h00}, /* 0x9b09 */
            {8'h00}, /* 0x9b08 */
            {8'h00}, /* 0x9b07 */
            {8'h00}, /* 0x9b06 */
            {8'h00}, /* 0x9b05 */
            {8'h00}, /* 0x9b04 */
            {8'h00}, /* 0x9b03 */
            {8'h00}, /* 0x9b02 */
            {8'h00}, /* 0x9b01 */
            {8'h00}, /* 0x9b00 */
            {8'h00}, /* 0x9aff */
            {8'h00}, /* 0x9afe */
            {8'h00}, /* 0x9afd */
            {8'h00}, /* 0x9afc */
            {8'h00}, /* 0x9afb */
            {8'h00}, /* 0x9afa */
            {8'h00}, /* 0x9af9 */
            {8'h00}, /* 0x9af8 */
            {8'h00}, /* 0x9af7 */
            {8'h00}, /* 0x9af6 */
            {8'h00}, /* 0x9af5 */
            {8'h00}, /* 0x9af4 */
            {8'h00}, /* 0x9af3 */
            {8'h00}, /* 0x9af2 */
            {8'h00}, /* 0x9af1 */
            {8'h00}, /* 0x9af0 */
            {8'h00}, /* 0x9aef */
            {8'h00}, /* 0x9aee */
            {8'h00}, /* 0x9aed */
            {8'h00}, /* 0x9aec */
            {8'h00}, /* 0x9aeb */
            {8'h00}, /* 0x9aea */
            {8'h00}, /* 0x9ae9 */
            {8'h00}, /* 0x9ae8 */
            {8'h00}, /* 0x9ae7 */
            {8'h00}, /* 0x9ae6 */
            {8'h00}, /* 0x9ae5 */
            {8'h00}, /* 0x9ae4 */
            {8'h00}, /* 0x9ae3 */
            {8'h00}, /* 0x9ae2 */
            {8'h00}, /* 0x9ae1 */
            {8'h00}, /* 0x9ae0 */
            {8'h00}, /* 0x9adf */
            {8'h00}, /* 0x9ade */
            {8'h00}, /* 0x9add */
            {8'h00}, /* 0x9adc */
            {8'h00}, /* 0x9adb */
            {8'h00}, /* 0x9ada */
            {8'h00}, /* 0x9ad9 */
            {8'h00}, /* 0x9ad8 */
            {8'h00}, /* 0x9ad7 */
            {8'h00}, /* 0x9ad6 */
            {8'h00}, /* 0x9ad5 */
            {8'h00}, /* 0x9ad4 */
            {8'h00}, /* 0x9ad3 */
            {8'h00}, /* 0x9ad2 */
            {8'h00}, /* 0x9ad1 */
            {8'h00}, /* 0x9ad0 */
            {8'h00}, /* 0x9acf */
            {8'h00}, /* 0x9ace */
            {8'h00}, /* 0x9acd */
            {8'h00}, /* 0x9acc */
            {8'h00}, /* 0x9acb */
            {8'h00}, /* 0x9aca */
            {8'h00}, /* 0x9ac9 */
            {8'h00}, /* 0x9ac8 */
            {8'h00}, /* 0x9ac7 */
            {8'h00}, /* 0x9ac6 */
            {8'h00}, /* 0x9ac5 */
            {8'h00}, /* 0x9ac4 */
            {8'h00}, /* 0x9ac3 */
            {8'h00}, /* 0x9ac2 */
            {8'h00}, /* 0x9ac1 */
            {8'h00}, /* 0x9ac0 */
            {8'h00}, /* 0x9abf */
            {8'h00}, /* 0x9abe */
            {8'h00}, /* 0x9abd */
            {8'h00}, /* 0x9abc */
            {8'h00}, /* 0x9abb */
            {8'h00}, /* 0x9aba */
            {8'h00}, /* 0x9ab9 */
            {8'h00}, /* 0x9ab8 */
            {8'h00}, /* 0x9ab7 */
            {8'h00}, /* 0x9ab6 */
            {8'h00}, /* 0x9ab5 */
            {8'h00}, /* 0x9ab4 */
            {8'h00}, /* 0x9ab3 */
            {8'h00}, /* 0x9ab2 */
            {8'h00}, /* 0x9ab1 */
            {8'h00}, /* 0x9ab0 */
            {8'h00}, /* 0x9aaf */
            {8'h00}, /* 0x9aae */
            {8'h00}, /* 0x9aad */
            {8'h00}, /* 0x9aac */
            {8'h00}, /* 0x9aab */
            {8'h00}, /* 0x9aaa */
            {8'h00}, /* 0x9aa9 */
            {8'h00}, /* 0x9aa8 */
            {8'h00}, /* 0x9aa7 */
            {8'h00}, /* 0x9aa6 */
            {8'h00}, /* 0x9aa5 */
            {8'h00}, /* 0x9aa4 */
            {8'h00}, /* 0x9aa3 */
            {8'h00}, /* 0x9aa2 */
            {8'h00}, /* 0x9aa1 */
            {8'h00}, /* 0x9aa0 */
            {8'h00}, /* 0x9a9f */
            {8'h00}, /* 0x9a9e */
            {8'h00}, /* 0x9a9d */
            {8'h00}, /* 0x9a9c */
            {8'h00}, /* 0x9a9b */
            {8'h00}, /* 0x9a9a */
            {8'h00}, /* 0x9a99 */
            {8'h00}, /* 0x9a98 */
            {8'h00}, /* 0x9a97 */
            {8'h00}, /* 0x9a96 */
            {8'h00}, /* 0x9a95 */
            {8'h00}, /* 0x9a94 */
            {8'h00}, /* 0x9a93 */
            {8'h00}, /* 0x9a92 */
            {8'h00}, /* 0x9a91 */
            {8'h00}, /* 0x9a90 */
            {8'h00}, /* 0x9a8f */
            {8'h00}, /* 0x9a8e */
            {8'h00}, /* 0x9a8d */
            {8'h00}, /* 0x9a8c */
            {8'h00}, /* 0x9a8b */
            {8'h00}, /* 0x9a8a */
            {8'h00}, /* 0x9a89 */
            {8'h00}, /* 0x9a88 */
            {8'h00}, /* 0x9a87 */
            {8'h00}, /* 0x9a86 */
            {8'h00}, /* 0x9a85 */
            {8'h00}, /* 0x9a84 */
            {8'h00}, /* 0x9a83 */
            {8'h00}, /* 0x9a82 */
            {8'h00}, /* 0x9a81 */
            {8'h00}, /* 0x9a80 */
            {8'h00}, /* 0x9a7f */
            {8'h00}, /* 0x9a7e */
            {8'h00}, /* 0x9a7d */
            {8'h00}, /* 0x9a7c */
            {8'h00}, /* 0x9a7b */
            {8'h00}, /* 0x9a7a */
            {8'h00}, /* 0x9a79 */
            {8'h00}, /* 0x9a78 */
            {8'h00}, /* 0x9a77 */
            {8'h00}, /* 0x9a76 */
            {8'h00}, /* 0x9a75 */
            {8'h00}, /* 0x9a74 */
            {8'h00}, /* 0x9a73 */
            {8'h00}, /* 0x9a72 */
            {8'h00}, /* 0x9a71 */
            {8'h00}, /* 0x9a70 */
            {8'h00}, /* 0x9a6f */
            {8'h00}, /* 0x9a6e */
            {8'h00}, /* 0x9a6d */
            {8'h00}, /* 0x9a6c */
            {8'h00}, /* 0x9a6b */
            {8'h00}, /* 0x9a6a */
            {8'h00}, /* 0x9a69 */
            {8'h00}, /* 0x9a68 */
            {8'h00}, /* 0x9a67 */
            {8'h00}, /* 0x9a66 */
            {8'h00}, /* 0x9a65 */
            {8'h00}, /* 0x9a64 */
            {8'h00}, /* 0x9a63 */
            {8'h00}, /* 0x9a62 */
            {8'h00}, /* 0x9a61 */
            {8'h00}, /* 0x9a60 */
            {8'h00}, /* 0x9a5f */
            {8'h00}, /* 0x9a5e */
            {8'h00}, /* 0x9a5d */
            {8'h00}, /* 0x9a5c */
            {8'h00}, /* 0x9a5b */
            {8'h00}, /* 0x9a5a */
            {8'h00}, /* 0x9a59 */
            {8'h00}, /* 0x9a58 */
            {8'h00}, /* 0x9a57 */
            {8'h00}, /* 0x9a56 */
            {8'h00}, /* 0x9a55 */
            {8'h00}, /* 0x9a54 */
            {8'h00}, /* 0x9a53 */
            {8'h00}, /* 0x9a52 */
            {8'h00}, /* 0x9a51 */
            {8'h00}, /* 0x9a50 */
            {8'h00}, /* 0x9a4f */
            {8'h00}, /* 0x9a4e */
            {8'h00}, /* 0x9a4d */
            {8'h00}, /* 0x9a4c */
            {8'h00}, /* 0x9a4b */
            {8'h00}, /* 0x9a4a */
            {8'h00}, /* 0x9a49 */
            {8'h00}, /* 0x9a48 */
            {8'h00}, /* 0x9a47 */
            {8'h00}, /* 0x9a46 */
            {8'h00}, /* 0x9a45 */
            {8'h00}, /* 0x9a44 */
            {8'h00}, /* 0x9a43 */
            {8'h00}, /* 0x9a42 */
            {8'h00}, /* 0x9a41 */
            {8'h00}, /* 0x9a40 */
            {8'h00}, /* 0x9a3f */
            {8'h00}, /* 0x9a3e */
            {8'h00}, /* 0x9a3d */
            {8'h00}, /* 0x9a3c */
            {8'h00}, /* 0x9a3b */
            {8'h00}, /* 0x9a3a */
            {8'h00}, /* 0x9a39 */
            {8'h00}, /* 0x9a38 */
            {8'h00}, /* 0x9a37 */
            {8'h00}, /* 0x9a36 */
            {8'h00}, /* 0x9a35 */
            {8'h00}, /* 0x9a34 */
            {8'h00}, /* 0x9a33 */
            {8'h00}, /* 0x9a32 */
            {8'h00}, /* 0x9a31 */
            {8'h00}, /* 0x9a30 */
            {8'h00}, /* 0x9a2f */
            {8'h00}, /* 0x9a2e */
            {8'h00}, /* 0x9a2d */
            {8'h00}, /* 0x9a2c */
            {8'h00}, /* 0x9a2b */
            {8'h00}, /* 0x9a2a */
            {8'h00}, /* 0x9a29 */
            {8'h00}, /* 0x9a28 */
            {8'h00}, /* 0x9a27 */
            {8'h00}, /* 0x9a26 */
            {8'h00}, /* 0x9a25 */
            {8'h00}, /* 0x9a24 */
            {8'h00}, /* 0x9a23 */
            {8'h00}, /* 0x9a22 */
            {8'h00}, /* 0x9a21 */
            {8'h00}, /* 0x9a20 */
            {8'h00}, /* 0x9a1f */
            {8'h00}, /* 0x9a1e */
            {8'h00}, /* 0x9a1d */
            {8'h00}, /* 0x9a1c */
            {8'h00}, /* 0x9a1b */
            {8'h00}, /* 0x9a1a */
            {8'h00}, /* 0x9a19 */
            {8'h00}, /* 0x9a18 */
            {8'h00}, /* 0x9a17 */
            {8'h00}, /* 0x9a16 */
            {8'h00}, /* 0x9a15 */
            {8'h00}, /* 0x9a14 */
            {8'h00}, /* 0x9a13 */
            {8'h00}, /* 0x9a12 */
            {8'h00}, /* 0x9a11 */
            {8'h00}, /* 0x9a10 */
            {8'h00}, /* 0x9a0f */
            {8'h00}, /* 0x9a0e */
            {8'h00}, /* 0x9a0d */
            {8'h00}, /* 0x9a0c */
            {8'h00}, /* 0x9a0b */
            {8'h00}, /* 0x9a0a */
            {8'h00}, /* 0x9a09 */
            {8'h00}, /* 0x9a08 */
            {8'h00}, /* 0x9a07 */
            {8'h00}, /* 0x9a06 */
            {8'h00}, /* 0x9a05 */
            {8'h00}, /* 0x9a04 */
            {8'h00}, /* 0x9a03 */
            {8'h00}, /* 0x9a02 */
            {8'h00}, /* 0x9a01 */
            {8'h00}, /* 0x9a00 */
            {8'h00}, /* 0x99ff */
            {8'h00}, /* 0x99fe */
            {8'h00}, /* 0x99fd */
            {8'h00}, /* 0x99fc */
            {8'h00}, /* 0x99fb */
            {8'h00}, /* 0x99fa */
            {8'h00}, /* 0x99f9 */
            {8'h00}, /* 0x99f8 */
            {8'h00}, /* 0x99f7 */
            {8'h00}, /* 0x99f6 */
            {8'h00}, /* 0x99f5 */
            {8'h00}, /* 0x99f4 */
            {8'h00}, /* 0x99f3 */
            {8'h00}, /* 0x99f2 */
            {8'h00}, /* 0x99f1 */
            {8'h00}, /* 0x99f0 */
            {8'h00}, /* 0x99ef */
            {8'h00}, /* 0x99ee */
            {8'h00}, /* 0x99ed */
            {8'h00}, /* 0x99ec */
            {8'h00}, /* 0x99eb */
            {8'h00}, /* 0x99ea */
            {8'h00}, /* 0x99e9 */
            {8'h00}, /* 0x99e8 */
            {8'h00}, /* 0x99e7 */
            {8'h00}, /* 0x99e6 */
            {8'h00}, /* 0x99e5 */
            {8'h00}, /* 0x99e4 */
            {8'h00}, /* 0x99e3 */
            {8'h00}, /* 0x99e2 */
            {8'h00}, /* 0x99e1 */
            {8'h00}, /* 0x99e0 */
            {8'h00}, /* 0x99df */
            {8'h00}, /* 0x99de */
            {8'h00}, /* 0x99dd */
            {8'h00}, /* 0x99dc */
            {8'h00}, /* 0x99db */
            {8'h00}, /* 0x99da */
            {8'h00}, /* 0x99d9 */
            {8'h00}, /* 0x99d8 */
            {8'h00}, /* 0x99d7 */
            {8'h00}, /* 0x99d6 */
            {8'h00}, /* 0x99d5 */
            {8'h00}, /* 0x99d4 */
            {8'h00}, /* 0x99d3 */
            {8'h00}, /* 0x99d2 */
            {8'h00}, /* 0x99d1 */
            {8'h00}, /* 0x99d0 */
            {8'h00}, /* 0x99cf */
            {8'h00}, /* 0x99ce */
            {8'h00}, /* 0x99cd */
            {8'h00}, /* 0x99cc */
            {8'h00}, /* 0x99cb */
            {8'h00}, /* 0x99ca */
            {8'h00}, /* 0x99c9 */
            {8'h00}, /* 0x99c8 */
            {8'h00}, /* 0x99c7 */
            {8'h00}, /* 0x99c6 */
            {8'h00}, /* 0x99c5 */
            {8'h00}, /* 0x99c4 */
            {8'h00}, /* 0x99c3 */
            {8'h00}, /* 0x99c2 */
            {8'h00}, /* 0x99c1 */
            {8'h00}, /* 0x99c0 */
            {8'h00}, /* 0x99bf */
            {8'h00}, /* 0x99be */
            {8'h00}, /* 0x99bd */
            {8'h00}, /* 0x99bc */
            {8'h00}, /* 0x99bb */
            {8'h00}, /* 0x99ba */
            {8'h00}, /* 0x99b9 */
            {8'h00}, /* 0x99b8 */
            {8'h00}, /* 0x99b7 */
            {8'h00}, /* 0x99b6 */
            {8'h00}, /* 0x99b5 */
            {8'h00}, /* 0x99b4 */
            {8'h00}, /* 0x99b3 */
            {8'h00}, /* 0x99b2 */
            {8'h00}, /* 0x99b1 */
            {8'h00}, /* 0x99b0 */
            {8'h00}, /* 0x99af */
            {8'h00}, /* 0x99ae */
            {8'h00}, /* 0x99ad */
            {8'h00}, /* 0x99ac */
            {8'h00}, /* 0x99ab */
            {8'h00}, /* 0x99aa */
            {8'h00}, /* 0x99a9 */
            {8'h00}, /* 0x99a8 */
            {8'h00}, /* 0x99a7 */
            {8'h00}, /* 0x99a6 */
            {8'h00}, /* 0x99a5 */
            {8'h00}, /* 0x99a4 */
            {8'h00}, /* 0x99a3 */
            {8'h00}, /* 0x99a2 */
            {8'h00}, /* 0x99a1 */
            {8'h00}, /* 0x99a0 */
            {8'h00}, /* 0x999f */
            {8'h00}, /* 0x999e */
            {8'h00}, /* 0x999d */
            {8'h00}, /* 0x999c */
            {8'h00}, /* 0x999b */
            {8'h00}, /* 0x999a */
            {8'h00}, /* 0x9999 */
            {8'h00}, /* 0x9998 */
            {8'h00}, /* 0x9997 */
            {8'h00}, /* 0x9996 */
            {8'h00}, /* 0x9995 */
            {8'h00}, /* 0x9994 */
            {8'h00}, /* 0x9993 */
            {8'h00}, /* 0x9992 */
            {8'h00}, /* 0x9991 */
            {8'h00}, /* 0x9990 */
            {8'h00}, /* 0x998f */
            {8'h00}, /* 0x998e */
            {8'h00}, /* 0x998d */
            {8'h00}, /* 0x998c */
            {8'h00}, /* 0x998b */
            {8'h00}, /* 0x998a */
            {8'h00}, /* 0x9989 */
            {8'h00}, /* 0x9988 */
            {8'h00}, /* 0x9987 */
            {8'h00}, /* 0x9986 */
            {8'h00}, /* 0x9985 */
            {8'h00}, /* 0x9984 */
            {8'h00}, /* 0x9983 */
            {8'h00}, /* 0x9982 */
            {8'h00}, /* 0x9981 */
            {8'h00}, /* 0x9980 */
            {8'h00}, /* 0x997f */
            {8'h00}, /* 0x997e */
            {8'h00}, /* 0x997d */
            {8'h00}, /* 0x997c */
            {8'h00}, /* 0x997b */
            {8'h00}, /* 0x997a */
            {8'h00}, /* 0x9979 */
            {8'h00}, /* 0x9978 */
            {8'h00}, /* 0x9977 */
            {8'h00}, /* 0x9976 */
            {8'h00}, /* 0x9975 */
            {8'h00}, /* 0x9974 */
            {8'h00}, /* 0x9973 */
            {8'h00}, /* 0x9972 */
            {8'h00}, /* 0x9971 */
            {8'h00}, /* 0x9970 */
            {8'h00}, /* 0x996f */
            {8'h00}, /* 0x996e */
            {8'h00}, /* 0x996d */
            {8'h00}, /* 0x996c */
            {8'h00}, /* 0x996b */
            {8'h00}, /* 0x996a */
            {8'h00}, /* 0x9969 */
            {8'h00}, /* 0x9968 */
            {8'h00}, /* 0x9967 */
            {8'h00}, /* 0x9966 */
            {8'h00}, /* 0x9965 */
            {8'h00}, /* 0x9964 */
            {8'h00}, /* 0x9963 */
            {8'h00}, /* 0x9962 */
            {8'h00}, /* 0x9961 */
            {8'h00}, /* 0x9960 */
            {8'h00}, /* 0x995f */
            {8'h00}, /* 0x995e */
            {8'h00}, /* 0x995d */
            {8'h00}, /* 0x995c */
            {8'h00}, /* 0x995b */
            {8'h00}, /* 0x995a */
            {8'h00}, /* 0x9959 */
            {8'h00}, /* 0x9958 */
            {8'h00}, /* 0x9957 */
            {8'h00}, /* 0x9956 */
            {8'h00}, /* 0x9955 */
            {8'h00}, /* 0x9954 */
            {8'h00}, /* 0x9953 */
            {8'h00}, /* 0x9952 */
            {8'h00}, /* 0x9951 */
            {8'h00}, /* 0x9950 */
            {8'h00}, /* 0x994f */
            {8'h00}, /* 0x994e */
            {8'h00}, /* 0x994d */
            {8'h00}, /* 0x994c */
            {8'h00}, /* 0x994b */
            {8'h00}, /* 0x994a */
            {8'h00}, /* 0x9949 */
            {8'h00}, /* 0x9948 */
            {8'h00}, /* 0x9947 */
            {8'h00}, /* 0x9946 */
            {8'h00}, /* 0x9945 */
            {8'h00}, /* 0x9944 */
            {8'h00}, /* 0x9943 */
            {8'h00}, /* 0x9942 */
            {8'h00}, /* 0x9941 */
            {8'h00}, /* 0x9940 */
            {8'h00}, /* 0x993f */
            {8'h00}, /* 0x993e */
            {8'h00}, /* 0x993d */
            {8'h00}, /* 0x993c */
            {8'h00}, /* 0x993b */
            {8'h00}, /* 0x993a */
            {8'h00}, /* 0x9939 */
            {8'h00}, /* 0x9938 */
            {8'h00}, /* 0x9937 */
            {8'h00}, /* 0x9936 */
            {8'h00}, /* 0x9935 */
            {8'h00}, /* 0x9934 */
            {8'h00}, /* 0x9933 */
            {8'h00}, /* 0x9932 */
            {8'h00}, /* 0x9931 */
            {8'h00}, /* 0x9930 */
            {8'h00}, /* 0x992f */
            {8'h00}, /* 0x992e */
            {8'h00}, /* 0x992d */
            {8'h00}, /* 0x992c */
            {8'h00}, /* 0x992b */
            {8'h00}, /* 0x992a */
            {8'h00}, /* 0x9929 */
            {8'h00}, /* 0x9928 */
            {8'h00}, /* 0x9927 */
            {8'h00}, /* 0x9926 */
            {8'h00}, /* 0x9925 */
            {8'h00}, /* 0x9924 */
            {8'h00}, /* 0x9923 */
            {8'h00}, /* 0x9922 */
            {8'h00}, /* 0x9921 */
            {8'h00}, /* 0x9920 */
            {8'h00}, /* 0x991f */
            {8'h00}, /* 0x991e */
            {8'h00}, /* 0x991d */
            {8'h00}, /* 0x991c */
            {8'h00}, /* 0x991b */
            {8'h00}, /* 0x991a */
            {8'h00}, /* 0x9919 */
            {8'h00}, /* 0x9918 */
            {8'h00}, /* 0x9917 */
            {8'h00}, /* 0x9916 */
            {8'h00}, /* 0x9915 */
            {8'h00}, /* 0x9914 */
            {8'h00}, /* 0x9913 */
            {8'h00}, /* 0x9912 */
            {8'h00}, /* 0x9911 */
            {8'h00}, /* 0x9910 */
            {8'h00}, /* 0x990f */
            {8'h00}, /* 0x990e */
            {8'h00}, /* 0x990d */
            {8'h00}, /* 0x990c */
            {8'h00}, /* 0x990b */
            {8'h00}, /* 0x990a */
            {8'h00}, /* 0x9909 */
            {8'h00}, /* 0x9908 */
            {8'h00}, /* 0x9907 */
            {8'h00}, /* 0x9906 */
            {8'h00}, /* 0x9905 */
            {8'h00}, /* 0x9904 */
            {8'h00}, /* 0x9903 */
            {8'h00}, /* 0x9902 */
            {8'h00}, /* 0x9901 */
            {8'h00}, /* 0x9900 */
            {8'h00}, /* 0x98ff */
            {8'h00}, /* 0x98fe */
            {8'h00}, /* 0x98fd */
            {8'h00}, /* 0x98fc */
            {8'h00}, /* 0x98fb */
            {8'h00}, /* 0x98fa */
            {8'h00}, /* 0x98f9 */
            {8'h00}, /* 0x98f8 */
            {8'h00}, /* 0x98f7 */
            {8'h00}, /* 0x98f6 */
            {8'h00}, /* 0x98f5 */
            {8'h00}, /* 0x98f4 */
            {8'h00}, /* 0x98f3 */
            {8'h00}, /* 0x98f2 */
            {8'h00}, /* 0x98f1 */
            {8'h00}, /* 0x98f0 */
            {8'h00}, /* 0x98ef */
            {8'h00}, /* 0x98ee */
            {8'h00}, /* 0x98ed */
            {8'h00}, /* 0x98ec */
            {8'h00}, /* 0x98eb */
            {8'h00}, /* 0x98ea */
            {8'h00}, /* 0x98e9 */
            {8'h00}, /* 0x98e8 */
            {8'h00}, /* 0x98e7 */
            {8'h00}, /* 0x98e6 */
            {8'h00}, /* 0x98e5 */
            {8'h00}, /* 0x98e4 */
            {8'h00}, /* 0x98e3 */
            {8'h00}, /* 0x98e2 */
            {8'h00}, /* 0x98e1 */
            {8'h00}, /* 0x98e0 */
            {8'h00}, /* 0x98df */
            {8'h00}, /* 0x98de */
            {8'h00}, /* 0x98dd */
            {8'h00}, /* 0x98dc */
            {8'h00}, /* 0x98db */
            {8'h00}, /* 0x98da */
            {8'h00}, /* 0x98d9 */
            {8'h00}, /* 0x98d8 */
            {8'h00}, /* 0x98d7 */
            {8'h00}, /* 0x98d6 */
            {8'h00}, /* 0x98d5 */
            {8'h00}, /* 0x98d4 */
            {8'h00}, /* 0x98d3 */
            {8'h00}, /* 0x98d2 */
            {8'h00}, /* 0x98d1 */
            {8'h00}, /* 0x98d0 */
            {8'h00}, /* 0x98cf */
            {8'h00}, /* 0x98ce */
            {8'h00}, /* 0x98cd */
            {8'h00}, /* 0x98cc */
            {8'h00}, /* 0x98cb */
            {8'h00}, /* 0x98ca */
            {8'h00}, /* 0x98c9 */
            {8'h00}, /* 0x98c8 */
            {8'h00}, /* 0x98c7 */
            {8'h00}, /* 0x98c6 */
            {8'h00}, /* 0x98c5 */
            {8'h00}, /* 0x98c4 */
            {8'h00}, /* 0x98c3 */
            {8'h00}, /* 0x98c2 */
            {8'h00}, /* 0x98c1 */
            {8'h00}, /* 0x98c0 */
            {8'h00}, /* 0x98bf */
            {8'h00}, /* 0x98be */
            {8'h00}, /* 0x98bd */
            {8'h00}, /* 0x98bc */
            {8'h00}, /* 0x98bb */
            {8'h00}, /* 0x98ba */
            {8'h00}, /* 0x98b9 */
            {8'h00}, /* 0x98b8 */
            {8'h00}, /* 0x98b7 */
            {8'h00}, /* 0x98b6 */
            {8'h00}, /* 0x98b5 */
            {8'h00}, /* 0x98b4 */
            {8'h00}, /* 0x98b3 */
            {8'h00}, /* 0x98b2 */
            {8'h00}, /* 0x98b1 */
            {8'h00}, /* 0x98b0 */
            {8'h00}, /* 0x98af */
            {8'h00}, /* 0x98ae */
            {8'h00}, /* 0x98ad */
            {8'h00}, /* 0x98ac */
            {8'h00}, /* 0x98ab */
            {8'h00}, /* 0x98aa */
            {8'h00}, /* 0x98a9 */
            {8'h00}, /* 0x98a8 */
            {8'h00}, /* 0x98a7 */
            {8'h00}, /* 0x98a6 */
            {8'h00}, /* 0x98a5 */
            {8'h00}, /* 0x98a4 */
            {8'h00}, /* 0x98a3 */
            {8'h00}, /* 0x98a2 */
            {8'h00}, /* 0x98a1 */
            {8'h00}, /* 0x98a0 */
            {8'h00}, /* 0x989f */
            {8'h00}, /* 0x989e */
            {8'h00}, /* 0x989d */
            {8'h00}, /* 0x989c */
            {8'h00}, /* 0x989b */
            {8'h00}, /* 0x989a */
            {8'h00}, /* 0x9899 */
            {8'h00}, /* 0x9898 */
            {8'h00}, /* 0x9897 */
            {8'h00}, /* 0x9896 */
            {8'h00}, /* 0x9895 */
            {8'h00}, /* 0x9894 */
            {8'h00}, /* 0x9893 */
            {8'h00}, /* 0x9892 */
            {8'h00}, /* 0x9891 */
            {8'h00}, /* 0x9890 */
            {8'h00}, /* 0x988f */
            {8'h00}, /* 0x988e */
            {8'h00}, /* 0x988d */
            {8'h00}, /* 0x988c */
            {8'h00}, /* 0x988b */
            {8'h00}, /* 0x988a */
            {8'h00}, /* 0x9889 */
            {8'h00}, /* 0x9888 */
            {8'h00}, /* 0x9887 */
            {8'h00}, /* 0x9886 */
            {8'h00}, /* 0x9885 */
            {8'h00}, /* 0x9884 */
            {8'h00}, /* 0x9883 */
            {8'h00}, /* 0x9882 */
            {8'h00}, /* 0x9881 */
            {8'h00}, /* 0x9880 */
            {8'h00}, /* 0x987f */
            {8'h00}, /* 0x987e */
            {8'h00}, /* 0x987d */
            {8'h00}, /* 0x987c */
            {8'h00}, /* 0x987b */
            {8'h00}, /* 0x987a */
            {8'h00}, /* 0x9879 */
            {8'h00}, /* 0x9878 */
            {8'h00}, /* 0x9877 */
            {8'h00}, /* 0x9876 */
            {8'h00}, /* 0x9875 */
            {8'h00}, /* 0x9874 */
            {8'h00}, /* 0x9873 */
            {8'h00}, /* 0x9872 */
            {8'h00}, /* 0x9871 */
            {8'h00}, /* 0x9870 */
            {8'h00}, /* 0x986f */
            {8'h00}, /* 0x986e */
            {8'h00}, /* 0x986d */
            {8'h00}, /* 0x986c */
            {8'h00}, /* 0x986b */
            {8'h00}, /* 0x986a */
            {8'h00}, /* 0x9869 */
            {8'h00}, /* 0x9868 */
            {8'h00}, /* 0x9867 */
            {8'h00}, /* 0x9866 */
            {8'h00}, /* 0x9865 */
            {8'h00}, /* 0x9864 */
            {8'h00}, /* 0x9863 */
            {8'h00}, /* 0x9862 */
            {8'h00}, /* 0x9861 */
            {8'h00}, /* 0x9860 */
            {8'h00}, /* 0x985f */
            {8'h00}, /* 0x985e */
            {8'h00}, /* 0x985d */
            {8'h00}, /* 0x985c */
            {8'h00}, /* 0x985b */
            {8'h00}, /* 0x985a */
            {8'h00}, /* 0x9859 */
            {8'h00}, /* 0x9858 */
            {8'h00}, /* 0x9857 */
            {8'h00}, /* 0x9856 */
            {8'h00}, /* 0x9855 */
            {8'h00}, /* 0x9854 */
            {8'h00}, /* 0x9853 */
            {8'h00}, /* 0x9852 */
            {8'h00}, /* 0x9851 */
            {8'h00}, /* 0x9850 */
            {8'h00}, /* 0x984f */
            {8'h00}, /* 0x984e */
            {8'h00}, /* 0x984d */
            {8'h00}, /* 0x984c */
            {8'h00}, /* 0x984b */
            {8'h00}, /* 0x984a */
            {8'h00}, /* 0x9849 */
            {8'h00}, /* 0x9848 */
            {8'h00}, /* 0x9847 */
            {8'h00}, /* 0x9846 */
            {8'h00}, /* 0x9845 */
            {8'h00}, /* 0x9844 */
            {8'h00}, /* 0x9843 */
            {8'h00}, /* 0x9842 */
            {8'h00}, /* 0x9841 */
            {8'h00}, /* 0x9840 */
            {8'h00}, /* 0x983f */
            {8'h00}, /* 0x983e */
            {8'h00}, /* 0x983d */
            {8'h00}, /* 0x983c */
            {8'h00}, /* 0x983b */
            {8'h00}, /* 0x983a */
            {8'h00}, /* 0x9839 */
            {8'h00}, /* 0x9838 */
            {8'h00}, /* 0x9837 */
            {8'h00}, /* 0x9836 */
            {8'h00}, /* 0x9835 */
            {8'h00}, /* 0x9834 */
            {8'h00}, /* 0x9833 */
            {8'h00}, /* 0x9832 */
            {8'h00}, /* 0x9831 */
            {8'h00}, /* 0x9830 */
            {8'h00}, /* 0x982f */
            {8'h00}, /* 0x982e */
            {8'h00}, /* 0x982d */
            {8'h00}, /* 0x982c */
            {8'h00}, /* 0x982b */
            {8'h00}, /* 0x982a */
            {8'h00}, /* 0x9829 */
            {8'h00}, /* 0x9828 */
            {8'h00}, /* 0x9827 */
            {8'h00}, /* 0x9826 */
            {8'h00}, /* 0x9825 */
            {8'h00}, /* 0x9824 */
            {8'h00}, /* 0x9823 */
            {8'h00}, /* 0x9822 */
            {8'h00}, /* 0x9821 */
            {8'h00}, /* 0x9820 */
            {8'h00}, /* 0x981f */
            {8'h00}, /* 0x981e */
            {8'h00}, /* 0x981d */
            {8'h00}, /* 0x981c */
            {8'h00}, /* 0x981b */
            {8'h00}, /* 0x981a */
            {8'h00}, /* 0x9819 */
            {8'h00}, /* 0x9818 */
            {8'h00}, /* 0x9817 */
            {8'h00}, /* 0x9816 */
            {8'h00}, /* 0x9815 */
            {8'h00}, /* 0x9814 */
            {8'h00}, /* 0x9813 */
            {8'h00}, /* 0x9812 */
            {8'h00}, /* 0x9811 */
            {8'h00}, /* 0x9810 */
            {8'h00}, /* 0x980f */
            {8'h00}, /* 0x980e */
            {8'h00}, /* 0x980d */
            {8'h00}, /* 0x980c */
            {8'h00}, /* 0x980b */
            {8'h00}, /* 0x980a */
            {8'h00}, /* 0x9809 */
            {8'h00}, /* 0x9808 */
            {8'h00}, /* 0x9807 */
            {8'h00}, /* 0x9806 */
            {8'h00}, /* 0x9805 */
            {8'h00}, /* 0x9804 */
            {8'h00}, /* 0x9803 */
            {8'h00}, /* 0x9802 */
            {8'h00}, /* 0x9801 */
            {8'h00}, /* 0x9800 */
            {8'h00}, /* 0x97ff */
            {8'h00}, /* 0x97fe */
            {8'h00}, /* 0x97fd */
            {8'h00}, /* 0x97fc */
            {8'h00}, /* 0x97fb */
            {8'h00}, /* 0x97fa */
            {8'h00}, /* 0x97f9 */
            {8'h00}, /* 0x97f8 */
            {8'h00}, /* 0x97f7 */
            {8'h00}, /* 0x97f6 */
            {8'h00}, /* 0x97f5 */
            {8'h00}, /* 0x97f4 */
            {8'h00}, /* 0x97f3 */
            {8'h00}, /* 0x97f2 */
            {8'h00}, /* 0x97f1 */
            {8'h00}, /* 0x97f0 */
            {8'h00}, /* 0x97ef */
            {8'h00}, /* 0x97ee */
            {8'h00}, /* 0x97ed */
            {8'h00}, /* 0x97ec */
            {8'h00}, /* 0x97eb */
            {8'h00}, /* 0x97ea */
            {8'h00}, /* 0x97e9 */
            {8'h00}, /* 0x97e8 */
            {8'h00}, /* 0x97e7 */
            {8'h00}, /* 0x97e6 */
            {8'h00}, /* 0x97e5 */
            {8'h00}, /* 0x97e4 */
            {8'h00}, /* 0x97e3 */
            {8'h00}, /* 0x97e2 */
            {8'h00}, /* 0x97e1 */
            {8'h00}, /* 0x97e0 */
            {8'h00}, /* 0x97df */
            {8'h00}, /* 0x97de */
            {8'h00}, /* 0x97dd */
            {8'h00}, /* 0x97dc */
            {8'h00}, /* 0x97db */
            {8'h00}, /* 0x97da */
            {8'h00}, /* 0x97d9 */
            {8'h00}, /* 0x97d8 */
            {8'h00}, /* 0x97d7 */
            {8'h00}, /* 0x97d6 */
            {8'h00}, /* 0x97d5 */
            {8'h00}, /* 0x97d4 */
            {8'h00}, /* 0x97d3 */
            {8'h00}, /* 0x97d2 */
            {8'h00}, /* 0x97d1 */
            {8'h00}, /* 0x97d0 */
            {8'h00}, /* 0x97cf */
            {8'h00}, /* 0x97ce */
            {8'h00}, /* 0x97cd */
            {8'h00}, /* 0x97cc */
            {8'h00}, /* 0x97cb */
            {8'h00}, /* 0x97ca */
            {8'h00}, /* 0x97c9 */
            {8'h00}, /* 0x97c8 */
            {8'h00}, /* 0x97c7 */
            {8'h00}, /* 0x97c6 */
            {8'h00}, /* 0x97c5 */
            {8'h00}, /* 0x97c4 */
            {8'h00}, /* 0x97c3 */
            {8'h00}, /* 0x97c2 */
            {8'h00}, /* 0x97c1 */
            {8'h00}, /* 0x97c0 */
            {8'h00}, /* 0x97bf */
            {8'h00}, /* 0x97be */
            {8'h00}, /* 0x97bd */
            {8'h00}, /* 0x97bc */
            {8'h00}, /* 0x97bb */
            {8'h00}, /* 0x97ba */
            {8'h00}, /* 0x97b9 */
            {8'h00}, /* 0x97b8 */
            {8'h00}, /* 0x97b7 */
            {8'h00}, /* 0x97b6 */
            {8'h00}, /* 0x97b5 */
            {8'h00}, /* 0x97b4 */
            {8'h00}, /* 0x97b3 */
            {8'h00}, /* 0x97b2 */
            {8'h00}, /* 0x97b1 */
            {8'h00}, /* 0x97b0 */
            {8'h00}, /* 0x97af */
            {8'h00}, /* 0x97ae */
            {8'h00}, /* 0x97ad */
            {8'h00}, /* 0x97ac */
            {8'h00}, /* 0x97ab */
            {8'h00}, /* 0x97aa */
            {8'h00}, /* 0x97a9 */
            {8'h00}, /* 0x97a8 */
            {8'h00}, /* 0x97a7 */
            {8'h00}, /* 0x97a6 */
            {8'h00}, /* 0x97a5 */
            {8'h00}, /* 0x97a4 */
            {8'h00}, /* 0x97a3 */
            {8'h00}, /* 0x97a2 */
            {8'h00}, /* 0x97a1 */
            {8'h00}, /* 0x97a0 */
            {8'h00}, /* 0x979f */
            {8'h00}, /* 0x979e */
            {8'h00}, /* 0x979d */
            {8'h00}, /* 0x979c */
            {8'h00}, /* 0x979b */
            {8'h00}, /* 0x979a */
            {8'h00}, /* 0x9799 */
            {8'h00}, /* 0x9798 */
            {8'h00}, /* 0x9797 */
            {8'h00}, /* 0x9796 */
            {8'h00}, /* 0x9795 */
            {8'h00}, /* 0x9794 */
            {8'h00}, /* 0x9793 */
            {8'h00}, /* 0x9792 */
            {8'h00}, /* 0x9791 */
            {8'h00}, /* 0x9790 */
            {8'h00}, /* 0x978f */
            {8'h00}, /* 0x978e */
            {8'h00}, /* 0x978d */
            {8'h00}, /* 0x978c */
            {8'h00}, /* 0x978b */
            {8'h00}, /* 0x978a */
            {8'h00}, /* 0x9789 */
            {8'h00}, /* 0x9788 */
            {8'h00}, /* 0x9787 */
            {8'h00}, /* 0x9786 */
            {8'h00}, /* 0x9785 */
            {8'h00}, /* 0x9784 */
            {8'h00}, /* 0x9783 */
            {8'h00}, /* 0x9782 */
            {8'h00}, /* 0x9781 */
            {8'h00}, /* 0x9780 */
            {8'h00}, /* 0x977f */
            {8'h00}, /* 0x977e */
            {8'h00}, /* 0x977d */
            {8'h00}, /* 0x977c */
            {8'h00}, /* 0x977b */
            {8'h00}, /* 0x977a */
            {8'h00}, /* 0x9779 */
            {8'h00}, /* 0x9778 */
            {8'h00}, /* 0x9777 */
            {8'h00}, /* 0x9776 */
            {8'h00}, /* 0x9775 */
            {8'h00}, /* 0x9774 */
            {8'h00}, /* 0x9773 */
            {8'h00}, /* 0x9772 */
            {8'h00}, /* 0x9771 */
            {8'h00}, /* 0x9770 */
            {8'h00}, /* 0x976f */
            {8'h00}, /* 0x976e */
            {8'h00}, /* 0x976d */
            {8'h00}, /* 0x976c */
            {8'h00}, /* 0x976b */
            {8'h00}, /* 0x976a */
            {8'h00}, /* 0x9769 */
            {8'h00}, /* 0x9768 */
            {8'h00}, /* 0x9767 */
            {8'h00}, /* 0x9766 */
            {8'h00}, /* 0x9765 */
            {8'h00}, /* 0x9764 */
            {8'h00}, /* 0x9763 */
            {8'h00}, /* 0x9762 */
            {8'h00}, /* 0x9761 */
            {8'h00}, /* 0x9760 */
            {8'h00}, /* 0x975f */
            {8'h00}, /* 0x975e */
            {8'h00}, /* 0x975d */
            {8'h00}, /* 0x975c */
            {8'h00}, /* 0x975b */
            {8'h00}, /* 0x975a */
            {8'h00}, /* 0x9759 */
            {8'h00}, /* 0x9758 */
            {8'h00}, /* 0x9757 */
            {8'h00}, /* 0x9756 */
            {8'h00}, /* 0x9755 */
            {8'h00}, /* 0x9754 */
            {8'h00}, /* 0x9753 */
            {8'h00}, /* 0x9752 */
            {8'h00}, /* 0x9751 */
            {8'h00}, /* 0x9750 */
            {8'h00}, /* 0x974f */
            {8'h00}, /* 0x974e */
            {8'h00}, /* 0x974d */
            {8'h00}, /* 0x974c */
            {8'h00}, /* 0x974b */
            {8'h00}, /* 0x974a */
            {8'h00}, /* 0x9749 */
            {8'h00}, /* 0x9748 */
            {8'h00}, /* 0x9747 */
            {8'h00}, /* 0x9746 */
            {8'h00}, /* 0x9745 */
            {8'h00}, /* 0x9744 */
            {8'h00}, /* 0x9743 */
            {8'h00}, /* 0x9742 */
            {8'h00}, /* 0x9741 */
            {8'h00}, /* 0x9740 */
            {8'h00}, /* 0x973f */
            {8'h00}, /* 0x973e */
            {8'h00}, /* 0x973d */
            {8'h00}, /* 0x973c */
            {8'h00}, /* 0x973b */
            {8'h00}, /* 0x973a */
            {8'h00}, /* 0x9739 */
            {8'h00}, /* 0x9738 */
            {8'h00}, /* 0x9737 */
            {8'h00}, /* 0x9736 */
            {8'h00}, /* 0x9735 */
            {8'h00}, /* 0x9734 */
            {8'h00}, /* 0x9733 */
            {8'h00}, /* 0x9732 */
            {8'h00}, /* 0x9731 */
            {8'h00}, /* 0x9730 */
            {8'h00}, /* 0x972f */
            {8'h00}, /* 0x972e */
            {8'h00}, /* 0x972d */
            {8'h00}, /* 0x972c */
            {8'h00}, /* 0x972b */
            {8'h00}, /* 0x972a */
            {8'h00}, /* 0x9729 */
            {8'h00}, /* 0x9728 */
            {8'h00}, /* 0x9727 */
            {8'h00}, /* 0x9726 */
            {8'h00}, /* 0x9725 */
            {8'h00}, /* 0x9724 */
            {8'h00}, /* 0x9723 */
            {8'h00}, /* 0x9722 */
            {8'h00}, /* 0x9721 */
            {8'h00}, /* 0x9720 */
            {8'h00}, /* 0x971f */
            {8'h00}, /* 0x971e */
            {8'h00}, /* 0x971d */
            {8'h00}, /* 0x971c */
            {8'h00}, /* 0x971b */
            {8'h00}, /* 0x971a */
            {8'h00}, /* 0x9719 */
            {8'h00}, /* 0x9718 */
            {8'h00}, /* 0x9717 */
            {8'h00}, /* 0x9716 */
            {8'h00}, /* 0x9715 */
            {8'h00}, /* 0x9714 */
            {8'h00}, /* 0x9713 */
            {8'h00}, /* 0x9712 */
            {8'h00}, /* 0x9711 */
            {8'h00}, /* 0x9710 */
            {8'h00}, /* 0x970f */
            {8'h00}, /* 0x970e */
            {8'h00}, /* 0x970d */
            {8'h00}, /* 0x970c */
            {8'h00}, /* 0x970b */
            {8'h00}, /* 0x970a */
            {8'h00}, /* 0x9709 */
            {8'h00}, /* 0x9708 */
            {8'h00}, /* 0x9707 */
            {8'h00}, /* 0x9706 */
            {8'h00}, /* 0x9705 */
            {8'h00}, /* 0x9704 */
            {8'h00}, /* 0x9703 */
            {8'h00}, /* 0x9702 */
            {8'h00}, /* 0x9701 */
            {8'h00}, /* 0x9700 */
            {8'h00}, /* 0x96ff */
            {8'h00}, /* 0x96fe */
            {8'h00}, /* 0x96fd */
            {8'h00}, /* 0x96fc */
            {8'h00}, /* 0x96fb */
            {8'h00}, /* 0x96fa */
            {8'h00}, /* 0x96f9 */
            {8'h00}, /* 0x96f8 */
            {8'h00}, /* 0x96f7 */
            {8'h00}, /* 0x96f6 */
            {8'h00}, /* 0x96f5 */
            {8'h00}, /* 0x96f4 */
            {8'h00}, /* 0x96f3 */
            {8'h00}, /* 0x96f2 */
            {8'h00}, /* 0x96f1 */
            {8'h00}, /* 0x96f0 */
            {8'h00}, /* 0x96ef */
            {8'h00}, /* 0x96ee */
            {8'h00}, /* 0x96ed */
            {8'h00}, /* 0x96ec */
            {8'h00}, /* 0x96eb */
            {8'h00}, /* 0x96ea */
            {8'h00}, /* 0x96e9 */
            {8'h00}, /* 0x96e8 */
            {8'h00}, /* 0x96e7 */
            {8'h00}, /* 0x96e6 */
            {8'h00}, /* 0x96e5 */
            {8'h00}, /* 0x96e4 */
            {8'h00}, /* 0x96e3 */
            {8'h00}, /* 0x96e2 */
            {8'h00}, /* 0x96e1 */
            {8'h00}, /* 0x96e0 */
            {8'h00}, /* 0x96df */
            {8'h00}, /* 0x96de */
            {8'h00}, /* 0x96dd */
            {8'h00}, /* 0x96dc */
            {8'h00}, /* 0x96db */
            {8'h00}, /* 0x96da */
            {8'h00}, /* 0x96d9 */
            {8'h00}, /* 0x96d8 */
            {8'h00}, /* 0x96d7 */
            {8'h00}, /* 0x96d6 */
            {8'h00}, /* 0x96d5 */
            {8'h00}, /* 0x96d4 */
            {8'h00}, /* 0x96d3 */
            {8'h00}, /* 0x96d2 */
            {8'h00}, /* 0x96d1 */
            {8'h00}, /* 0x96d0 */
            {8'h00}, /* 0x96cf */
            {8'h00}, /* 0x96ce */
            {8'h00}, /* 0x96cd */
            {8'h00}, /* 0x96cc */
            {8'h00}, /* 0x96cb */
            {8'h00}, /* 0x96ca */
            {8'h00}, /* 0x96c9 */
            {8'h00}, /* 0x96c8 */
            {8'h00}, /* 0x96c7 */
            {8'h00}, /* 0x96c6 */
            {8'h00}, /* 0x96c5 */
            {8'h00}, /* 0x96c4 */
            {8'h00}, /* 0x96c3 */
            {8'h00}, /* 0x96c2 */
            {8'h00}, /* 0x96c1 */
            {8'h00}, /* 0x96c0 */
            {8'h00}, /* 0x96bf */
            {8'h00}, /* 0x96be */
            {8'h00}, /* 0x96bd */
            {8'h00}, /* 0x96bc */
            {8'h00}, /* 0x96bb */
            {8'h00}, /* 0x96ba */
            {8'h00}, /* 0x96b9 */
            {8'h00}, /* 0x96b8 */
            {8'h00}, /* 0x96b7 */
            {8'h00}, /* 0x96b6 */
            {8'h00}, /* 0x96b5 */
            {8'h00}, /* 0x96b4 */
            {8'h00}, /* 0x96b3 */
            {8'h00}, /* 0x96b2 */
            {8'h00}, /* 0x96b1 */
            {8'h00}, /* 0x96b0 */
            {8'h00}, /* 0x96af */
            {8'h00}, /* 0x96ae */
            {8'h00}, /* 0x96ad */
            {8'h00}, /* 0x96ac */
            {8'h00}, /* 0x96ab */
            {8'h00}, /* 0x96aa */
            {8'h00}, /* 0x96a9 */
            {8'h00}, /* 0x96a8 */
            {8'h00}, /* 0x96a7 */
            {8'h00}, /* 0x96a6 */
            {8'h00}, /* 0x96a5 */
            {8'h00}, /* 0x96a4 */
            {8'h00}, /* 0x96a3 */
            {8'h00}, /* 0x96a2 */
            {8'h00}, /* 0x96a1 */
            {8'h00}, /* 0x96a0 */
            {8'h00}, /* 0x969f */
            {8'h00}, /* 0x969e */
            {8'h00}, /* 0x969d */
            {8'h00}, /* 0x969c */
            {8'h00}, /* 0x969b */
            {8'h00}, /* 0x969a */
            {8'h00}, /* 0x9699 */
            {8'h00}, /* 0x9698 */
            {8'h00}, /* 0x9697 */
            {8'h00}, /* 0x9696 */
            {8'h00}, /* 0x9695 */
            {8'h00}, /* 0x9694 */
            {8'h00}, /* 0x9693 */
            {8'h00}, /* 0x9692 */
            {8'h00}, /* 0x9691 */
            {8'h00}, /* 0x9690 */
            {8'h00}, /* 0x968f */
            {8'h00}, /* 0x968e */
            {8'h00}, /* 0x968d */
            {8'h00}, /* 0x968c */
            {8'h00}, /* 0x968b */
            {8'h00}, /* 0x968a */
            {8'h00}, /* 0x9689 */
            {8'h00}, /* 0x9688 */
            {8'h00}, /* 0x9687 */
            {8'h00}, /* 0x9686 */
            {8'h00}, /* 0x9685 */
            {8'h00}, /* 0x9684 */
            {8'h00}, /* 0x9683 */
            {8'h00}, /* 0x9682 */
            {8'h00}, /* 0x9681 */
            {8'h00}, /* 0x9680 */
            {8'h00}, /* 0x967f */
            {8'h00}, /* 0x967e */
            {8'h00}, /* 0x967d */
            {8'h00}, /* 0x967c */
            {8'h00}, /* 0x967b */
            {8'h00}, /* 0x967a */
            {8'h00}, /* 0x9679 */
            {8'h00}, /* 0x9678 */
            {8'h00}, /* 0x9677 */
            {8'h00}, /* 0x9676 */
            {8'h00}, /* 0x9675 */
            {8'h00}, /* 0x9674 */
            {8'h00}, /* 0x9673 */
            {8'h00}, /* 0x9672 */
            {8'h00}, /* 0x9671 */
            {8'h00}, /* 0x9670 */
            {8'h00}, /* 0x966f */
            {8'h00}, /* 0x966e */
            {8'h00}, /* 0x966d */
            {8'h00}, /* 0x966c */
            {8'h00}, /* 0x966b */
            {8'h00}, /* 0x966a */
            {8'h00}, /* 0x9669 */
            {8'h00}, /* 0x9668 */
            {8'h00}, /* 0x9667 */
            {8'h00}, /* 0x9666 */
            {8'h00}, /* 0x9665 */
            {8'h00}, /* 0x9664 */
            {8'h00}, /* 0x9663 */
            {8'h00}, /* 0x9662 */
            {8'h00}, /* 0x9661 */
            {8'h00}, /* 0x9660 */
            {8'h00}, /* 0x965f */
            {8'h00}, /* 0x965e */
            {8'h00}, /* 0x965d */
            {8'h00}, /* 0x965c */
            {8'h00}, /* 0x965b */
            {8'h00}, /* 0x965a */
            {8'h00}, /* 0x9659 */
            {8'h00}, /* 0x9658 */
            {8'h00}, /* 0x9657 */
            {8'h00}, /* 0x9656 */
            {8'h00}, /* 0x9655 */
            {8'h00}, /* 0x9654 */
            {8'h00}, /* 0x9653 */
            {8'h00}, /* 0x9652 */
            {8'h00}, /* 0x9651 */
            {8'h00}, /* 0x9650 */
            {8'h00}, /* 0x964f */
            {8'h00}, /* 0x964e */
            {8'h00}, /* 0x964d */
            {8'h00}, /* 0x964c */
            {8'h00}, /* 0x964b */
            {8'h00}, /* 0x964a */
            {8'h00}, /* 0x9649 */
            {8'h00}, /* 0x9648 */
            {8'h00}, /* 0x9647 */
            {8'h00}, /* 0x9646 */
            {8'h00}, /* 0x9645 */
            {8'h00}, /* 0x9644 */
            {8'h00}, /* 0x9643 */
            {8'h00}, /* 0x9642 */
            {8'h00}, /* 0x9641 */
            {8'h00}, /* 0x9640 */
            {8'h00}, /* 0x963f */
            {8'h00}, /* 0x963e */
            {8'h00}, /* 0x963d */
            {8'h00}, /* 0x963c */
            {8'h00}, /* 0x963b */
            {8'h00}, /* 0x963a */
            {8'h00}, /* 0x9639 */
            {8'h00}, /* 0x9638 */
            {8'h00}, /* 0x9637 */
            {8'h00}, /* 0x9636 */
            {8'h00}, /* 0x9635 */
            {8'h00}, /* 0x9634 */
            {8'h00}, /* 0x9633 */
            {8'h00}, /* 0x9632 */
            {8'h00}, /* 0x9631 */
            {8'h00}, /* 0x9630 */
            {8'h00}, /* 0x962f */
            {8'h00}, /* 0x962e */
            {8'h00}, /* 0x962d */
            {8'h00}, /* 0x962c */
            {8'h00}, /* 0x962b */
            {8'h00}, /* 0x962a */
            {8'h00}, /* 0x9629 */
            {8'h00}, /* 0x9628 */
            {8'h00}, /* 0x9627 */
            {8'h00}, /* 0x9626 */
            {8'h00}, /* 0x9625 */
            {8'h00}, /* 0x9624 */
            {8'h00}, /* 0x9623 */
            {8'h00}, /* 0x9622 */
            {8'h00}, /* 0x9621 */
            {8'h00}, /* 0x9620 */
            {8'h00}, /* 0x961f */
            {8'h00}, /* 0x961e */
            {8'h00}, /* 0x961d */
            {8'h00}, /* 0x961c */
            {8'h00}, /* 0x961b */
            {8'h00}, /* 0x961a */
            {8'h00}, /* 0x9619 */
            {8'h00}, /* 0x9618 */
            {8'h00}, /* 0x9617 */
            {8'h00}, /* 0x9616 */
            {8'h00}, /* 0x9615 */
            {8'h00}, /* 0x9614 */
            {8'h00}, /* 0x9613 */
            {8'h00}, /* 0x9612 */
            {8'h00}, /* 0x9611 */
            {8'h00}, /* 0x9610 */
            {8'h00}, /* 0x960f */
            {8'h00}, /* 0x960e */
            {8'h00}, /* 0x960d */
            {8'h00}, /* 0x960c */
            {8'h00}, /* 0x960b */
            {8'h00}, /* 0x960a */
            {8'h00}, /* 0x9609 */
            {8'h00}, /* 0x9608 */
            {8'h00}, /* 0x9607 */
            {8'h00}, /* 0x9606 */
            {8'h00}, /* 0x9605 */
            {8'h00}, /* 0x9604 */
            {8'h00}, /* 0x9603 */
            {8'h00}, /* 0x9602 */
            {8'h00}, /* 0x9601 */
            {8'h00}, /* 0x9600 */
            {8'h00}, /* 0x95ff */
            {8'h00}, /* 0x95fe */
            {8'h00}, /* 0x95fd */
            {8'h00}, /* 0x95fc */
            {8'h00}, /* 0x95fb */
            {8'h00}, /* 0x95fa */
            {8'h00}, /* 0x95f9 */
            {8'h00}, /* 0x95f8 */
            {8'h00}, /* 0x95f7 */
            {8'h00}, /* 0x95f6 */
            {8'h00}, /* 0x95f5 */
            {8'h00}, /* 0x95f4 */
            {8'h00}, /* 0x95f3 */
            {8'h00}, /* 0x95f2 */
            {8'h00}, /* 0x95f1 */
            {8'h00}, /* 0x95f0 */
            {8'h00}, /* 0x95ef */
            {8'h00}, /* 0x95ee */
            {8'h00}, /* 0x95ed */
            {8'h00}, /* 0x95ec */
            {8'h00}, /* 0x95eb */
            {8'h00}, /* 0x95ea */
            {8'h00}, /* 0x95e9 */
            {8'h00}, /* 0x95e8 */
            {8'h00}, /* 0x95e7 */
            {8'h00}, /* 0x95e6 */
            {8'h00}, /* 0x95e5 */
            {8'h00}, /* 0x95e4 */
            {8'h00}, /* 0x95e3 */
            {8'h00}, /* 0x95e2 */
            {8'h00}, /* 0x95e1 */
            {8'h00}, /* 0x95e0 */
            {8'h00}, /* 0x95df */
            {8'h00}, /* 0x95de */
            {8'h00}, /* 0x95dd */
            {8'h00}, /* 0x95dc */
            {8'h00}, /* 0x95db */
            {8'h00}, /* 0x95da */
            {8'h00}, /* 0x95d9 */
            {8'h00}, /* 0x95d8 */
            {8'h00}, /* 0x95d7 */
            {8'h00}, /* 0x95d6 */
            {8'h00}, /* 0x95d5 */
            {8'h00}, /* 0x95d4 */
            {8'h00}, /* 0x95d3 */
            {8'h00}, /* 0x95d2 */
            {8'h00}, /* 0x95d1 */
            {8'h00}, /* 0x95d0 */
            {8'h00}, /* 0x95cf */
            {8'h00}, /* 0x95ce */
            {8'h00}, /* 0x95cd */
            {8'h00}, /* 0x95cc */
            {8'h00}, /* 0x95cb */
            {8'h00}, /* 0x95ca */
            {8'h00}, /* 0x95c9 */
            {8'h00}, /* 0x95c8 */
            {8'h00}, /* 0x95c7 */
            {8'h00}, /* 0x95c6 */
            {8'h00}, /* 0x95c5 */
            {8'h00}, /* 0x95c4 */
            {8'h00}, /* 0x95c3 */
            {8'h00}, /* 0x95c2 */
            {8'h00}, /* 0x95c1 */
            {8'h00}, /* 0x95c0 */
            {8'h00}, /* 0x95bf */
            {8'h00}, /* 0x95be */
            {8'h00}, /* 0x95bd */
            {8'h00}, /* 0x95bc */
            {8'h00}, /* 0x95bb */
            {8'h00}, /* 0x95ba */
            {8'h00}, /* 0x95b9 */
            {8'h00}, /* 0x95b8 */
            {8'h00}, /* 0x95b7 */
            {8'h00}, /* 0x95b6 */
            {8'h00}, /* 0x95b5 */
            {8'h00}, /* 0x95b4 */
            {8'h00}, /* 0x95b3 */
            {8'h00}, /* 0x95b2 */
            {8'h00}, /* 0x95b1 */
            {8'h00}, /* 0x95b0 */
            {8'h00}, /* 0x95af */
            {8'h00}, /* 0x95ae */
            {8'h00}, /* 0x95ad */
            {8'h00}, /* 0x95ac */
            {8'h00}, /* 0x95ab */
            {8'h00}, /* 0x95aa */
            {8'h00}, /* 0x95a9 */
            {8'h00}, /* 0x95a8 */
            {8'h00}, /* 0x95a7 */
            {8'h00}, /* 0x95a6 */
            {8'h00}, /* 0x95a5 */
            {8'h00}, /* 0x95a4 */
            {8'h00}, /* 0x95a3 */
            {8'h00}, /* 0x95a2 */
            {8'h00}, /* 0x95a1 */
            {8'h00}, /* 0x95a0 */
            {8'h00}, /* 0x959f */
            {8'h00}, /* 0x959e */
            {8'h00}, /* 0x959d */
            {8'h00}, /* 0x959c */
            {8'h00}, /* 0x959b */
            {8'h00}, /* 0x959a */
            {8'h00}, /* 0x9599 */
            {8'h00}, /* 0x9598 */
            {8'h00}, /* 0x9597 */
            {8'h00}, /* 0x9596 */
            {8'h00}, /* 0x9595 */
            {8'h00}, /* 0x9594 */
            {8'h00}, /* 0x9593 */
            {8'h00}, /* 0x9592 */
            {8'h00}, /* 0x9591 */
            {8'h00}, /* 0x9590 */
            {8'h00}, /* 0x958f */
            {8'h00}, /* 0x958e */
            {8'h00}, /* 0x958d */
            {8'h00}, /* 0x958c */
            {8'h00}, /* 0x958b */
            {8'h00}, /* 0x958a */
            {8'h00}, /* 0x9589 */
            {8'h00}, /* 0x9588 */
            {8'h00}, /* 0x9587 */
            {8'h00}, /* 0x9586 */
            {8'h00}, /* 0x9585 */
            {8'h00}, /* 0x9584 */
            {8'h00}, /* 0x9583 */
            {8'h00}, /* 0x9582 */
            {8'h00}, /* 0x9581 */
            {8'h00}, /* 0x9580 */
            {8'h00}, /* 0x957f */
            {8'h00}, /* 0x957e */
            {8'h00}, /* 0x957d */
            {8'h00}, /* 0x957c */
            {8'h00}, /* 0x957b */
            {8'h00}, /* 0x957a */
            {8'h00}, /* 0x9579 */
            {8'h00}, /* 0x9578 */
            {8'h00}, /* 0x9577 */
            {8'h00}, /* 0x9576 */
            {8'h00}, /* 0x9575 */
            {8'h00}, /* 0x9574 */
            {8'h00}, /* 0x9573 */
            {8'h00}, /* 0x9572 */
            {8'h00}, /* 0x9571 */
            {8'h00}, /* 0x9570 */
            {8'h00}, /* 0x956f */
            {8'h00}, /* 0x956e */
            {8'h00}, /* 0x956d */
            {8'h00}, /* 0x956c */
            {8'h00}, /* 0x956b */
            {8'h00}, /* 0x956a */
            {8'h00}, /* 0x9569 */
            {8'h00}, /* 0x9568 */
            {8'h00}, /* 0x9567 */
            {8'h00}, /* 0x9566 */
            {8'h00}, /* 0x9565 */
            {8'h00}, /* 0x9564 */
            {8'h00}, /* 0x9563 */
            {8'h00}, /* 0x9562 */
            {8'h00}, /* 0x9561 */
            {8'h00}, /* 0x9560 */
            {8'h00}, /* 0x955f */
            {8'h00}, /* 0x955e */
            {8'h00}, /* 0x955d */
            {8'h00}, /* 0x955c */
            {8'h00}, /* 0x955b */
            {8'h00}, /* 0x955a */
            {8'h00}, /* 0x9559 */
            {8'h00}, /* 0x9558 */
            {8'h00}, /* 0x9557 */
            {8'h00}, /* 0x9556 */
            {8'h00}, /* 0x9555 */
            {8'h00}, /* 0x9554 */
            {8'h00}, /* 0x9553 */
            {8'h00}, /* 0x9552 */
            {8'h00}, /* 0x9551 */
            {8'h00}, /* 0x9550 */
            {8'h00}, /* 0x954f */
            {8'h00}, /* 0x954e */
            {8'h00}, /* 0x954d */
            {8'h00}, /* 0x954c */
            {8'h00}, /* 0x954b */
            {8'h00}, /* 0x954a */
            {8'h00}, /* 0x9549 */
            {8'h00}, /* 0x9548 */
            {8'h00}, /* 0x9547 */
            {8'h00}, /* 0x9546 */
            {8'h00}, /* 0x9545 */
            {8'h00}, /* 0x9544 */
            {8'h00}, /* 0x9543 */
            {8'h00}, /* 0x9542 */
            {8'h00}, /* 0x9541 */
            {8'h00}, /* 0x9540 */
            {8'h00}, /* 0x953f */
            {8'h00}, /* 0x953e */
            {8'h00}, /* 0x953d */
            {8'h00}, /* 0x953c */
            {8'h00}, /* 0x953b */
            {8'h00}, /* 0x953a */
            {8'h00}, /* 0x9539 */
            {8'h00}, /* 0x9538 */
            {8'h00}, /* 0x9537 */
            {8'h00}, /* 0x9536 */
            {8'h00}, /* 0x9535 */
            {8'h00}, /* 0x9534 */
            {8'h00}, /* 0x9533 */
            {8'h00}, /* 0x9532 */
            {8'h00}, /* 0x9531 */
            {8'h00}, /* 0x9530 */
            {8'h00}, /* 0x952f */
            {8'h00}, /* 0x952e */
            {8'h00}, /* 0x952d */
            {8'h00}, /* 0x952c */
            {8'h00}, /* 0x952b */
            {8'h00}, /* 0x952a */
            {8'h00}, /* 0x9529 */
            {8'h00}, /* 0x9528 */
            {8'h00}, /* 0x9527 */
            {8'h00}, /* 0x9526 */
            {8'h00}, /* 0x9525 */
            {8'h00}, /* 0x9524 */
            {8'h00}, /* 0x9523 */
            {8'h00}, /* 0x9522 */
            {8'h00}, /* 0x9521 */
            {8'h00}, /* 0x9520 */
            {8'h00}, /* 0x951f */
            {8'h00}, /* 0x951e */
            {8'h00}, /* 0x951d */
            {8'h00}, /* 0x951c */
            {8'h00}, /* 0x951b */
            {8'h00}, /* 0x951a */
            {8'h00}, /* 0x9519 */
            {8'h00}, /* 0x9518 */
            {8'h00}, /* 0x9517 */
            {8'h00}, /* 0x9516 */
            {8'h00}, /* 0x9515 */
            {8'h00}, /* 0x9514 */
            {8'h00}, /* 0x9513 */
            {8'h00}, /* 0x9512 */
            {8'h00}, /* 0x9511 */
            {8'h00}, /* 0x9510 */
            {8'h00}, /* 0x950f */
            {8'h00}, /* 0x950e */
            {8'h00}, /* 0x950d */
            {8'h00}, /* 0x950c */
            {8'h00}, /* 0x950b */
            {8'h00}, /* 0x950a */
            {8'h00}, /* 0x9509 */
            {8'h00}, /* 0x9508 */
            {8'h00}, /* 0x9507 */
            {8'h00}, /* 0x9506 */
            {8'h00}, /* 0x9505 */
            {8'h00}, /* 0x9504 */
            {8'h00}, /* 0x9503 */
            {8'h00}, /* 0x9502 */
            {8'h00}, /* 0x9501 */
            {8'h00}, /* 0x9500 */
            {8'h00}, /* 0x94ff */
            {8'h00}, /* 0x94fe */
            {8'h00}, /* 0x94fd */
            {8'h00}, /* 0x94fc */
            {8'h00}, /* 0x94fb */
            {8'h00}, /* 0x94fa */
            {8'h00}, /* 0x94f9 */
            {8'h00}, /* 0x94f8 */
            {8'h00}, /* 0x94f7 */
            {8'h00}, /* 0x94f6 */
            {8'h00}, /* 0x94f5 */
            {8'h00}, /* 0x94f4 */
            {8'h00}, /* 0x94f3 */
            {8'h00}, /* 0x94f2 */
            {8'h00}, /* 0x94f1 */
            {8'h00}, /* 0x94f0 */
            {8'h00}, /* 0x94ef */
            {8'h00}, /* 0x94ee */
            {8'h00}, /* 0x94ed */
            {8'h00}, /* 0x94ec */
            {8'h00}, /* 0x94eb */
            {8'h00}, /* 0x94ea */
            {8'h00}, /* 0x94e9 */
            {8'h00}, /* 0x94e8 */
            {8'h00}, /* 0x94e7 */
            {8'h00}, /* 0x94e6 */
            {8'h00}, /* 0x94e5 */
            {8'h00}, /* 0x94e4 */
            {8'h00}, /* 0x94e3 */
            {8'h00}, /* 0x94e2 */
            {8'h00}, /* 0x94e1 */
            {8'h00}, /* 0x94e0 */
            {8'h00}, /* 0x94df */
            {8'h00}, /* 0x94de */
            {8'h00}, /* 0x94dd */
            {8'h00}, /* 0x94dc */
            {8'h00}, /* 0x94db */
            {8'h00}, /* 0x94da */
            {8'h00}, /* 0x94d9 */
            {8'h00}, /* 0x94d8 */
            {8'h00}, /* 0x94d7 */
            {8'h00}, /* 0x94d6 */
            {8'h00}, /* 0x94d5 */
            {8'h00}, /* 0x94d4 */
            {8'h00}, /* 0x94d3 */
            {8'h00}, /* 0x94d2 */
            {8'h00}, /* 0x94d1 */
            {8'h00}, /* 0x94d0 */
            {8'h00}, /* 0x94cf */
            {8'h00}, /* 0x94ce */
            {8'h00}, /* 0x94cd */
            {8'h00}, /* 0x94cc */
            {8'h00}, /* 0x94cb */
            {8'h00}, /* 0x94ca */
            {8'h00}, /* 0x94c9 */
            {8'h00}, /* 0x94c8 */
            {8'h00}, /* 0x94c7 */
            {8'h00}, /* 0x94c6 */
            {8'h00}, /* 0x94c5 */
            {8'h00}, /* 0x94c4 */
            {8'h00}, /* 0x94c3 */
            {8'h00}, /* 0x94c2 */
            {8'h00}, /* 0x94c1 */
            {8'h00}, /* 0x94c0 */
            {8'h00}, /* 0x94bf */
            {8'h00}, /* 0x94be */
            {8'h00}, /* 0x94bd */
            {8'h00}, /* 0x94bc */
            {8'h00}, /* 0x94bb */
            {8'h00}, /* 0x94ba */
            {8'h00}, /* 0x94b9 */
            {8'h00}, /* 0x94b8 */
            {8'h00}, /* 0x94b7 */
            {8'h00}, /* 0x94b6 */
            {8'h00}, /* 0x94b5 */
            {8'h00}, /* 0x94b4 */
            {8'h00}, /* 0x94b3 */
            {8'h00}, /* 0x94b2 */
            {8'h00}, /* 0x94b1 */
            {8'h00}, /* 0x94b0 */
            {8'h00}, /* 0x94af */
            {8'h00}, /* 0x94ae */
            {8'h00}, /* 0x94ad */
            {8'h00}, /* 0x94ac */
            {8'h00}, /* 0x94ab */
            {8'h00}, /* 0x94aa */
            {8'h00}, /* 0x94a9 */
            {8'h00}, /* 0x94a8 */
            {8'h00}, /* 0x94a7 */
            {8'h00}, /* 0x94a6 */
            {8'h00}, /* 0x94a5 */
            {8'h00}, /* 0x94a4 */
            {8'h00}, /* 0x94a3 */
            {8'h00}, /* 0x94a2 */
            {8'h00}, /* 0x94a1 */
            {8'h00}, /* 0x94a0 */
            {8'h00}, /* 0x949f */
            {8'h00}, /* 0x949e */
            {8'h00}, /* 0x949d */
            {8'h00}, /* 0x949c */
            {8'h00}, /* 0x949b */
            {8'h00}, /* 0x949a */
            {8'h00}, /* 0x9499 */
            {8'h00}, /* 0x9498 */
            {8'h00}, /* 0x9497 */
            {8'h00}, /* 0x9496 */
            {8'h00}, /* 0x9495 */
            {8'h00}, /* 0x9494 */
            {8'h00}, /* 0x9493 */
            {8'h00}, /* 0x9492 */
            {8'h00}, /* 0x9491 */
            {8'h00}, /* 0x9490 */
            {8'h00}, /* 0x948f */
            {8'h00}, /* 0x948e */
            {8'h00}, /* 0x948d */
            {8'h00}, /* 0x948c */
            {8'h00}, /* 0x948b */
            {8'h00}, /* 0x948a */
            {8'h00}, /* 0x9489 */
            {8'h00}, /* 0x9488 */
            {8'h00}, /* 0x9487 */
            {8'h00}, /* 0x9486 */
            {8'h00}, /* 0x9485 */
            {8'h00}, /* 0x9484 */
            {8'h00}, /* 0x9483 */
            {8'h00}, /* 0x9482 */
            {8'h00}, /* 0x9481 */
            {8'h00}, /* 0x9480 */
            {8'h00}, /* 0x947f */
            {8'h00}, /* 0x947e */
            {8'h00}, /* 0x947d */
            {8'h00}, /* 0x947c */
            {8'h00}, /* 0x947b */
            {8'h00}, /* 0x947a */
            {8'h00}, /* 0x9479 */
            {8'h00}, /* 0x9478 */
            {8'h00}, /* 0x9477 */
            {8'h00}, /* 0x9476 */
            {8'h00}, /* 0x9475 */
            {8'h00}, /* 0x9474 */
            {8'h00}, /* 0x9473 */
            {8'h00}, /* 0x9472 */
            {8'h00}, /* 0x9471 */
            {8'h00}, /* 0x9470 */
            {8'h00}, /* 0x946f */
            {8'h00}, /* 0x946e */
            {8'h00}, /* 0x946d */
            {8'h00}, /* 0x946c */
            {8'h00}, /* 0x946b */
            {8'h00}, /* 0x946a */
            {8'h00}, /* 0x9469 */
            {8'h00}, /* 0x9468 */
            {8'h00}, /* 0x9467 */
            {8'h00}, /* 0x9466 */
            {8'h00}, /* 0x9465 */
            {8'h00}, /* 0x9464 */
            {8'h00}, /* 0x9463 */
            {8'h00}, /* 0x9462 */
            {8'h00}, /* 0x9461 */
            {8'h00}, /* 0x9460 */
            {8'h00}, /* 0x945f */
            {8'h00}, /* 0x945e */
            {8'h00}, /* 0x945d */
            {8'h00}, /* 0x945c */
            {8'h00}, /* 0x945b */
            {8'h00}, /* 0x945a */
            {8'h00}, /* 0x9459 */
            {8'h00}, /* 0x9458 */
            {8'h00}, /* 0x9457 */
            {8'h00}, /* 0x9456 */
            {8'h00}, /* 0x9455 */
            {8'h00}, /* 0x9454 */
            {8'h00}, /* 0x9453 */
            {8'h00}, /* 0x9452 */
            {8'h00}, /* 0x9451 */
            {8'h00}, /* 0x9450 */
            {8'h00}, /* 0x944f */
            {8'h00}, /* 0x944e */
            {8'h00}, /* 0x944d */
            {8'h00}, /* 0x944c */
            {8'h00}, /* 0x944b */
            {8'h00}, /* 0x944a */
            {8'h00}, /* 0x9449 */
            {8'h00}, /* 0x9448 */
            {8'h00}, /* 0x9447 */
            {8'h00}, /* 0x9446 */
            {8'h00}, /* 0x9445 */
            {8'h00}, /* 0x9444 */
            {8'h00}, /* 0x9443 */
            {8'h00}, /* 0x9442 */
            {8'h00}, /* 0x9441 */
            {8'h00}, /* 0x9440 */
            {8'h00}, /* 0x943f */
            {8'h00}, /* 0x943e */
            {8'h00}, /* 0x943d */
            {8'h00}, /* 0x943c */
            {8'h00}, /* 0x943b */
            {8'h00}, /* 0x943a */
            {8'h00}, /* 0x9439 */
            {8'h00}, /* 0x9438 */
            {8'h00}, /* 0x9437 */
            {8'h00}, /* 0x9436 */
            {8'h00}, /* 0x9435 */
            {8'h00}, /* 0x9434 */
            {8'h00}, /* 0x9433 */
            {8'h00}, /* 0x9432 */
            {8'h00}, /* 0x9431 */
            {8'h00}, /* 0x9430 */
            {8'h00}, /* 0x942f */
            {8'h00}, /* 0x942e */
            {8'h00}, /* 0x942d */
            {8'h00}, /* 0x942c */
            {8'h00}, /* 0x942b */
            {8'h00}, /* 0x942a */
            {8'h00}, /* 0x9429 */
            {8'h00}, /* 0x9428 */
            {8'h00}, /* 0x9427 */
            {8'h00}, /* 0x9426 */
            {8'h00}, /* 0x9425 */
            {8'h00}, /* 0x9424 */
            {8'h00}, /* 0x9423 */
            {8'h00}, /* 0x9422 */
            {8'h00}, /* 0x9421 */
            {8'h00}, /* 0x9420 */
            {8'h00}, /* 0x941f */
            {8'h00}, /* 0x941e */
            {8'h00}, /* 0x941d */
            {8'h00}, /* 0x941c */
            {8'h00}, /* 0x941b */
            {8'h00}, /* 0x941a */
            {8'h00}, /* 0x9419 */
            {8'h00}, /* 0x9418 */
            {8'h00}, /* 0x9417 */
            {8'h00}, /* 0x9416 */
            {8'h00}, /* 0x9415 */
            {8'h00}, /* 0x9414 */
            {8'h00}, /* 0x9413 */
            {8'h00}, /* 0x9412 */
            {8'h00}, /* 0x9411 */
            {8'h00}, /* 0x9410 */
            {8'h00}, /* 0x940f */
            {8'h00}, /* 0x940e */
            {8'h00}, /* 0x940d */
            {8'h00}, /* 0x940c */
            {8'h00}, /* 0x940b */
            {8'h00}, /* 0x940a */
            {8'h00}, /* 0x9409 */
            {8'h00}, /* 0x9408 */
            {8'h00}, /* 0x9407 */
            {8'h00}, /* 0x9406 */
            {8'h00}, /* 0x9405 */
            {8'h00}, /* 0x9404 */
            {8'h00}, /* 0x9403 */
            {8'h00}, /* 0x9402 */
            {8'h00}, /* 0x9401 */
            {8'h00}, /* 0x9400 */
            {8'h00}, /* 0x93ff */
            {8'h00}, /* 0x93fe */
            {8'h00}, /* 0x93fd */
            {8'h00}, /* 0x93fc */
            {8'h00}, /* 0x93fb */
            {8'h00}, /* 0x93fa */
            {8'h00}, /* 0x93f9 */
            {8'h00}, /* 0x93f8 */
            {8'h00}, /* 0x93f7 */
            {8'h00}, /* 0x93f6 */
            {8'h00}, /* 0x93f5 */
            {8'h00}, /* 0x93f4 */
            {8'h00}, /* 0x93f3 */
            {8'h00}, /* 0x93f2 */
            {8'h00}, /* 0x93f1 */
            {8'h00}, /* 0x93f0 */
            {8'h00}, /* 0x93ef */
            {8'h00}, /* 0x93ee */
            {8'h00}, /* 0x93ed */
            {8'h00}, /* 0x93ec */
            {8'h00}, /* 0x93eb */
            {8'h00}, /* 0x93ea */
            {8'h00}, /* 0x93e9 */
            {8'h00}, /* 0x93e8 */
            {8'h00}, /* 0x93e7 */
            {8'h00}, /* 0x93e6 */
            {8'h00}, /* 0x93e5 */
            {8'h00}, /* 0x93e4 */
            {8'h00}, /* 0x93e3 */
            {8'h00}, /* 0x93e2 */
            {8'h00}, /* 0x93e1 */
            {8'h00}, /* 0x93e0 */
            {8'h00}, /* 0x93df */
            {8'h00}, /* 0x93de */
            {8'h00}, /* 0x93dd */
            {8'h00}, /* 0x93dc */
            {8'h00}, /* 0x93db */
            {8'h00}, /* 0x93da */
            {8'h00}, /* 0x93d9 */
            {8'h00}, /* 0x93d8 */
            {8'h00}, /* 0x93d7 */
            {8'h00}, /* 0x93d6 */
            {8'h00}, /* 0x93d5 */
            {8'h00}, /* 0x93d4 */
            {8'h00}, /* 0x93d3 */
            {8'h00}, /* 0x93d2 */
            {8'h00}, /* 0x93d1 */
            {8'h00}, /* 0x93d0 */
            {8'h00}, /* 0x93cf */
            {8'h00}, /* 0x93ce */
            {8'h00}, /* 0x93cd */
            {8'h00}, /* 0x93cc */
            {8'h00}, /* 0x93cb */
            {8'h00}, /* 0x93ca */
            {8'h00}, /* 0x93c9 */
            {8'h00}, /* 0x93c8 */
            {8'h00}, /* 0x93c7 */
            {8'h00}, /* 0x93c6 */
            {8'h00}, /* 0x93c5 */
            {8'h00}, /* 0x93c4 */
            {8'h00}, /* 0x93c3 */
            {8'h00}, /* 0x93c2 */
            {8'h00}, /* 0x93c1 */
            {8'h00}, /* 0x93c0 */
            {8'h00}, /* 0x93bf */
            {8'h00}, /* 0x93be */
            {8'h00}, /* 0x93bd */
            {8'h00}, /* 0x93bc */
            {8'h00}, /* 0x93bb */
            {8'h00}, /* 0x93ba */
            {8'h00}, /* 0x93b9 */
            {8'h00}, /* 0x93b8 */
            {8'h00}, /* 0x93b7 */
            {8'h00}, /* 0x93b6 */
            {8'h00}, /* 0x93b5 */
            {8'h00}, /* 0x93b4 */
            {8'h00}, /* 0x93b3 */
            {8'h00}, /* 0x93b2 */
            {8'h00}, /* 0x93b1 */
            {8'h00}, /* 0x93b0 */
            {8'h00}, /* 0x93af */
            {8'h00}, /* 0x93ae */
            {8'h00}, /* 0x93ad */
            {8'h00}, /* 0x93ac */
            {8'h00}, /* 0x93ab */
            {8'h00}, /* 0x93aa */
            {8'h00}, /* 0x93a9 */
            {8'h00}, /* 0x93a8 */
            {8'h00}, /* 0x93a7 */
            {8'h00}, /* 0x93a6 */
            {8'h00}, /* 0x93a5 */
            {8'h00}, /* 0x93a4 */
            {8'h00}, /* 0x93a3 */
            {8'h00}, /* 0x93a2 */
            {8'h00}, /* 0x93a1 */
            {8'h00}, /* 0x93a0 */
            {8'h00}, /* 0x939f */
            {8'h00}, /* 0x939e */
            {8'h00}, /* 0x939d */
            {8'h00}, /* 0x939c */
            {8'h00}, /* 0x939b */
            {8'h00}, /* 0x939a */
            {8'h00}, /* 0x9399 */
            {8'h00}, /* 0x9398 */
            {8'h00}, /* 0x9397 */
            {8'h00}, /* 0x9396 */
            {8'h00}, /* 0x9395 */
            {8'h00}, /* 0x9394 */
            {8'h00}, /* 0x9393 */
            {8'h00}, /* 0x9392 */
            {8'h00}, /* 0x9391 */
            {8'h00}, /* 0x9390 */
            {8'h00}, /* 0x938f */
            {8'h00}, /* 0x938e */
            {8'h00}, /* 0x938d */
            {8'h00}, /* 0x938c */
            {8'h00}, /* 0x938b */
            {8'h00}, /* 0x938a */
            {8'h00}, /* 0x9389 */
            {8'h00}, /* 0x9388 */
            {8'h00}, /* 0x9387 */
            {8'h00}, /* 0x9386 */
            {8'h00}, /* 0x9385 */
            {8'h00}, /* 0x9384 */
            {8'h00}, /* 0x9383 */
            {8'h00}, /* 0x9382 */
            {8'h00}, /* 0x9381 */
            {8'h00}, /* 0x9380 */
            {8'h00}, /* 0x937f */
            {8'h00}, /* 0x937e */
            {8'h00}, /* 0x937d */
            {8'h00}, /* 0x937c */
            {8'h00}, /* 0x937b */
            {8'h00}, /* 0x937a */
            {8'h00}, /* 0x9379 */
            {8'h00}, /* 0x9378 */
            {8'h00}, /* 0x9377 */
            {8'h00}, /* 0x9376 */
            {8'h00}, /* 0x9375 */
            {8'h00}, /* 0x9374 */
            {8'h00}, /* 0x9373 */
            {8'h00}, /* 0x9372 */
            {8'h00}, /* 0x9371 */
            {8'h00}, /* 0x9370 */
            {8'h00}, /* 0x936f */
            {8'h00}, /* 0x936e */
            {8'h00}, /* 0x936d */
            {8'h00}, /* 0x936c */
            {8'h00}, /* 0x936b */
            {8'h00}, /* 0x936a */
            {8'h00}, /* 0x9369 */
            {8'h00}, /* 0x9368 */
            {8'h00}, /* 0x9367 */
            {8'h00}, /* 0x9366 */
            {8'h00}, /* 0x9365 */
            {8'h00}, /* 0x9364 */
            {8'h00}, /* 0x9363 */
            {8'h00}, /* 0x9362 */
            {8'h00}, /* 0x9361 */
            {8'h00}, /* 0x9360 */
            {8'h00}, /* 0x935f */
            {8'h00}, /* 0x935e */
            {8'h00}, /* 0x935d */
            {8'h00}, /* 0x935c */
            {8'h00}, /* 0x935b */
            {8'h00}, /* 0x935a */
            {8'h00}, /* 0x9359 */
            {8'h00}, /* 0x9358 */
            {8'h00}, /* 0x9357 */
            {8'h00}, /* 0x9356 */
            {8'h00}, /* 0x9355 */
            {8'h00}, /* 0x9354 */
            {8'h00}, /* 0x9353 */
            {8'h00}, /* 0x9352 */
            {8'h00}, /* 0x9351 */
            {8'h00}, /* 0x9350 */
            {8'h00}, /* 0x934f */
            {8'h00}, /* 0x934e */
            {8'h00}, /* 0x934d */
            {8'h00}, /* 0x934c */
            {8'h00}, /* 0x934b */
            {8'h00}, /* 0x934a */
            {8'h00}, /* 0x9349 */
            {8'h00}, /* 0x9348 */
            {8'h00}, /* 0x9347 */
            {8'h00}, /* 0x9346 */
            {8'h00}, /* 0x9345 */
            {8'h00}, /* 0x9344 */
            {8'h00}, /* 0x9343 */
            {8'h00}, /* 0x9342 */
            {8'h00}, /* 0x9341 */
            {8'h00}, /* 0x9340 */
            {8'h00}, /* 0x933f */
            {8'h00}, /* 0x933e */
            {8'h00}, /* 0x933d */
            {8'h00}, /* 0x933c */
            {8'h00}, /* 0x933b */
            {8'h00}, /* 0x933a */
            {8'h00}, /* 0x9339 */
            {8'h00}, /* 0x9338 */
            {8'h00}, /* 0x9337 */
            {8'h00}, /* 0x9336 */
            {8'h00}, /* 0x9335 */
            {8'h00}, /* 0x9334 */
            {8'h00}, /* 0x9333 */
            {8'h00}, /* 0x9332 */
            {8'h00}, /* 0x9331 */
            {8'h00}, /* 0x9330 */
            {8'h00}, /* 0x932f */
            {8'h00}, /* 0x932e */
            {8'h00}, /* 0x932d */
            {8'h00}, /* 0x932c */
            {8'h00}, /* 0x932b */
            {8'h00}, /* 0x932a */
            {8'h00}, /* 0x9329 */
            {8'h00}, /* 0x9328 */
            {8'h00}, /* 0x9327 */
            {8'h00}, /* 0x9326 */
            {8'h00}, /* 0x9325 */
            {8'h00}, /* 0x9324 */
            {8'h00}, /* 0x9323 */
            {8'h00}, /* 0x9322 */
            {8'h00}, /* 0x9321 */
            {8'h00}, /* 0x9320 */
            {8'h00}, /* 0x931f */
            {8'h00}, /* 0x931e */
            {8'h00}, /* 0x931d */
            {8'h00}, /* 0x931c */
            {8'h00}, /* 0x931b */
            {8'h00}, /* 0x931a */
            {8'h00}, /* 0x9319 */
            {8'h00}, /* 0x9318 */
            {8'h00}, /* 0x9317 */
            {8'h00}, /* 0x9316 */
            {8'h00}, /* 0x9315 */
            {8'h00}, /* 0x9314 */
            {8'h00}, /* 0x9313 */
            {8'h00}, /* 0x9312 */
            {8'h00}, /* 0x9311 */
            {8'h00}, /* 0x9310 */
            {8'h00}, /* 0x930f */
            {8'h00}, /* 0x930e */
            {8'h00}, /* 0x930d */
            {8'h00}, /* 0x930c */
            {8'h00}, /* 0x930b */
            {8'h00}, /* 0x930a */
            {8'h00}, /* 0x9309 */
            {8'h00}, /* 0x9308 */
            {8'h00}, /* 0x9307 */
            {8'h00}, /* 0x9306 */
            {8'h00}, /* 0x9305 */
            {8'h00}, /* 0x9304 */
            {8'h00}, /* 0x9303 */
            {8'h00}, /* 0x9302 */
            {8'h00}, /* 0x9301 */
            {8'h00}, /* 0x9300 */
            {8'h00}, /* 0x92ff */
            {8'h00}, /* 0x92fe */
            {8'h00}, /* 0x92fd */
            {8'h00}, /* 0x92fc */
            {8'h00}, /* 0x92fb */
            {8'h00}, /* 0x92fa */
            {8'h00}, /* 0x92f9 */
            {8'h00}, /* 0x92f8 */
            {8'h00}, /* 0x92f7 */
            {8'h00}, /* 0x92f6 */
            {8'h00}, /* 0x92f5 */
            {8'h00}, /* 0x92f4 */
            {8'h00}, /* 0x92f3 */
            {8'h00}, /* 0x92f2 */
            {8'h00}, /* 0x92f1 */
            {8'h00}, /* 0x92f0 */
            {8'h00}, /* 0x92ef */
            {8'h00}, /* 0x92ee */
            {8'h00}, /* 0x92ed */
            {8'h00}, /* 0x92ec */
            {8'h00}, /* 0x92eb */
            {8'h00}, /* 0x92ea */
            {8'h00}, /* 0x92e9 */
            {8'h00}, /* 0x92e8 */
            {8'h00}, /* 0x92e7 */
            {8'h00}, /* 0x92e6 */
            {8'h00}, /* 0x92e5 */
            {8'h00}, /* 0x92e4 */
            {8'h00}, /* 0x92e3 */
            {8'h00}, /* 0x92e2 */
            {8'h00}, /* 0x92e1 */
            {8'h00}, /* 0x92e0 */
            {8'h00}, /* 0x92df */
            {8'h00}, /* 0x92de */
            {8'h00}, /* 0x92dd */
            {8'h00}, /* 0x92dc */
            {8'h00}, /* 0x92db */
            {8'h00}, /* 0x92da */
            {8'h00}, /* 0x92d9 */
            {8'h00}, /* 0x92d8 */
            {8'h00}, /* 0x92d7 */
            {8'h00}, /* 0x92d6 */
            {8'h00}, /* 0x92d5 */
            {8'h00}, /* 0x92d4 */
            {8'h00}, /* 0x92d3 */
            {8'h00}, /* 0x92d2 */
            {8'h00}, /* 0x92d1 */
            {8'h00}, /* 0x92d0 */
            {8'h00}, /* 0x92cf */
            {8'h00}, /* 0x92ce */
            {8'h00}, /* 0x92cd */
            {8'h00}, /* 0x92cc */
            {8'h00}, /* 0x92cb */
            {8'h00}, /* 0x92ca */
            {8'h00}, /* 0x92c9 */
            {8'h00}, /* 0x92c8 */
            {8'h00}, /* 0x92c7 */
            {8'h00}, /* 0x92c6 */
            {8'h00}, /* 0x92c5 */
            {8'h00}, /* 0x92c4 */
            {8'h00}, /* 0x92c3 */
            {8'h00}, /* 0x92c2 */
            {8'h00}, /* 0x92c1 */
            {8'h00}, /* 0x92c0 */
            {8'h00}, /* 0x92bf */
            {8'h00}, /* 0x92be */
            {8'h00}, /* 0x92bd */
            {8'h00}, /* 0x92bc */
            {8'h00}, /* 0x92bb */
            {8'h00}, /* 0x92ba */
            {8'h00}, /* 0x92b9 */
            {8'h00}, /* 0x92b8 */
            {8'h00}, /* 0x92b7 */
            {8'h00}, /* 0x92b6 */
            {8'h00}, /* 0x92b5 */
            {8'h00}, /* 0x92b4 */
            {8'h00}, /* 0x92b3 */
            {8'h00}, /* 0x92b2 */
            {8'h00}, /* 0x92b1 */
            {8'h00}, /* 0x92b0 */
            {8'h00}, /* 0x92af */
            {8'h00}, /* 0x92ae */
            {8'h00}, /* 0x92ad */
            {8'h00}, /* 0x92ac */
            {8'h00}, /* 0x92ab */
            {8'h00}, /* 0x92aa */
            {8'h00}, /* 0x92a9 */
            {8'h00}, /* 0x92a8 */
            {8'h00}, /* 0x92a7 */
            {8'h00}, /* 0x92a6 */
            {8'h00}, /* 0x92a5 */
            {8'h00}, /* 0x92a4 */
            {8'h00}, /* 0x92a3 */
            {8'h00}, /* 0x92a2 */
            {8'h00}, /* 0x92a1 */
            {8'h00}, /* 0x92a0 */
            {8'h00}, /* 0x929f */
            {8'h00}, /* 0x929e */
            {8'h00}, /* 0x929d */
            {8'h00}, /* 0x929c */
            {8'h00}, /* 0x929b */
            {8'h00}, /* 0x929a */
            {8'h00}, /* 0x9299 */
            {8'h00}, /* 0x9298 */
            {8'h00}, /* 0x9297 */
            {8'h00}, /* 0x9296 */
            {8'h00}, /* 0x9295 */
            {8'h00}, /* 0x9294 */
            {8'h00}, /* 0x9293 */
            {8'h00}, /* 0x9292 */
            {8'h00}, /* 0x9291 */
            {8'h00}, /* 0x9290 */
            {8'h00}, /* 0x928f */
            {8'h00}, /* 0x928e */
            {8'h00}, /* 0x928d */
            {8'h00}, /* 0x928c */
            {8'h00}, /* 0x928b */
            {8'h00}, /* 0x928a */
            {8'h00}, /* 0x9289 */
            {8'h00}, /* 0x9288 */
            {8'h00}, /* 0x9287 */
            {8'h00}, /* 0x9286 */
            {8'h00}, /* 0x9285 */
            {8'h00}, /* 0x9284 */
            {8'h00}, /* 0x9283 */
            {8'h00}, /* 0x9282 */
            {8'h00}, /* 0x9281 */
            {8'h00}, /* 0x9280 */
            {8'h00}, /* 0x927f */
            {8'h00}, /* 0x927e */
            {8'h00}, /* 0x927d */
            {8'h00}, /* 0x927c */
            {8'h00}, /* 0x927b */
            {8'h00}, /* 0x927a */
            {8'h00}, /* 0x9279 */
            {8'h00}, /* 0x9278 */
            {8'h00}, /* 0x9277 */
            {8'h00}, /* 0x9276 */
            {8'h00}, /* 0x9275 */
            {8'h00}, /* 0x9274 */
            {8'h00}, /* 0x9273 */
            {8'h00}, /* 0x9272 */
            {8'h00}, /* 0x9271 */
            {8'h00}, /* 0x9270 */
            {8'h00}, /* 0x926f */
            {8'h00}, /* 0x926e */
            {8'h00}, /* 0x926d */
            {8'h00}, /* 0x926c */
            {8'h00}, /* 0x926b */
            {8'h00}, /* 0x926a */
            {8'h00}, /* 0x9269 */
            {8'h00}, /* 0x9268 */
            {8'h00}, /* 0x9267 */
            {8'h00}, /* 0x9266 */
            {8'h00}, /* 0x9265 */
            {8'h00}, /* 0x9264 */
            {8'h00}, /* 0x9263 */
            {8'h00}, /* 0x9262 */
            {8'h00}, /* 0x9261 */
            {8'h00}, /* 0x9260 */
            {8'h00}, /* 0x925f */
            {8'h00}, /* 0x925e */
            {8'h00}, /* 0x925d */
            {8'h00}, /* 0x925c */
            {8'h00}, /* 0x925b */
            {8'h00}, /* 0x925a */
            {8'h00}, /* 0x9259 */
            {8'h00}, /* 0x9258 */
            {8'h00}, /* 0x9257 */
            {8'h00}, /* 0x9256 */
            {8'h00}, /* 0x9255 */
            {8'h00}, /* 0x9254 */
            {8'h00}, /* 0x9253 */
            {8'h00}, /* 0x9252 */
            {8'h00}, /* 0x9251 */
            {8'h00}, /* 0x9250 */
            {8'h00}, /* 0x924f */
            {8'h00}, /* 0x924e */
            {8'h00}, /* 0x924d */
            {8'h00}, /* 0x924c */
            {8'h00}, /* 0x924b */
            {8'h00}, /* 0x924a */
            {8'h00}, /* 0x9249 */
            {8'h00}, /* 0x9248 */
            {8'h00}, /* 0x9247 */
            {8'h00}, /* 0x9246 */
            {8'h00}, /* 0x9245 */
            {8'h00}, /* 0x9244 */
            {8'h00}, /* 0x9243 */
            {8'h00}, /* 0x9242 */
            {8'h00}, /* 0x9241 */
            {8'h00}, /* 0x9240 */
            {8'h00}, /* 0x923f */
            {8'h00}, /* 0x923e */
            {8'h00}, /* 0x923d */
            {8'h00}, /* 0x923c */
            {8'h00}, /* 0x923b */
            {8'h00}, /* 0x923a */
            {8'h00}, /* 0x9239 */
            {8'h00}, /* 0x9238 */
            {8'h00}, /* 0x9237 */
            {8'h00}, /* 0x9236 */
            {8'h00}, /* 0x9235 */
            {8'h00}, /* 0x9234 */
            {8'h00}, /* 0x9233 */
            {8'h00}, /* 0x9232 */
            {8'h00}, /* 0x9231 */
            {8'h00}, /* 0x9230 */
            {8'h00}, /* 0x922f */
            {8'h00}, /* 0x922e */
            {8'h00}, /* 0x922d */
            {8'h00}, /* 0x922c */
            {8'h00}, /* 0x922b */
            {8'h00}, /* 0x922a */
            {8'h00}, /* 0x9229 */
            {8'h00}, /* 0x9228 */
            {8'h00}, /* 0x9227 */
            {8'h00}, /* 0x9226 */
            {8'h00}, /* 0x9225 */
            {8'h00}, /* 0x9224 */
            {8'h00}, /* 0x9223 */
            {8'h00}, /* 0x9222 */
            {8'h00}, /* 0x9221 */
            {8'h00}, /* 0x9220 */
            {8'h00}, /* 0x921f */
            {8'h00}, /* 0x921e */
            {8'h00}, /* 0x921d */
            {8'h00}, /* 0x921c */
            {8'h00}, /* 0x921b */
            {8'h00}, /* 0x921a */
            {8'h00}, /* 0x9219 */
            {8'h00}, /* 0x9218 */
            {8'h00}, /* 0x9217 */
            {8'h00}, /* 0x9216 */
            {8'h00}, /* 0x9215 */
            {8'h00}, /* 0x9214 */
            {8'h00}, /* 0x9213 */
            {8'h00}, /* 0x9212 */
            {8'h00}, /* 0x9211 */
            {8'h00}, /* 0x9210 */
            {8'h00}, /* 0x920f */
            {8'h00}, /* 0x920e */
            {8'h00}, /* 0x920d */
            {8'h00}, /* 0x920c */
            {8'h00}, /* 0x920b */
            {8'h00}, /* 0x920a */
            {8'h00}, /* 0x9209 */
            {8'h00}, /* 0x9208 */
            {8'h00}, /* 0x9207 */
            {8'h00}, /* 0x9206 */
            {8'h00}, /* 0x9205 */
            {8'h00}, /* 0x9204 */
            {8'h00}, /* 0x9203 */
            {8'h00}, /* 0x9202 */
            {8'h00}, /* 0x9201 */
            {8'h00}, /* 0x9200 */
            {8'h00}, /* 0x91ff */
            {8'h00}, /* 0x91fe */
            {8'h00}, /* 0x91fd */
            {8'h00}, /* 0x91fc */
            {8'h00}, /* 0x91fb */
            {8'h00}, /* 0x91fa */
            {8'h00}, /* 0x91f9 */
            {8'h00}, /* 0x91f8 */
            {8'h00}, /* 0x91f7 */
            {8'h00}, /* 0x91f6 */
            {8'h00}, /* 0x91f5 */
            {8'h00}, /* 0x91f4 */
            {8'h00}, /* 0x91f3 */
            {8'h00}, /* 0x91f2 */
            {8'h00}, /* 0x91f1 */
            {8'h00}, /* 0x91f0 */
            {8'h00}, /* 0x91ef */
            {8'h00}, /* 0x91ee */
            {8'h00}, /* 0x91ed */
            {8'h00}, /* 0x91ec */
            {8'h00}, /* 0x91eb */
            {8'h00}, /* 0x91ea */
            {8'h00}, /* 0x91e9 */
            {8'h00}, /* 0x91e8 */
            {8'h00}, /* 0x91e7 */
            {8'h00}, /* 0x91e6 */
            {8'h00}, /* 0x91e5 */
            {8'h00}, /* 0x91e4 */
            {8'h00}, /* 0x91e3 */
            {8'h00}, /* 0x91e2 */
            {8'h00}, /* 0x91e1 */
            {8'h00}, /* 0x91e0 */
            {8'h00}, /* 0x91df */
            {8'h00}, /* 0x91de */
            {8'h00}, /* 0x91dd */
            {8'h00}, /* 0x91dc */
            {8'h00}, /* 0x91db */
            {8'h00}, /* 0x91da */
            {8'h00}, /* 0x91d9 */
            {8'h00}, /* 0x91d8 */
            {8'h00}, /* 0x91d7 */
            {8'h00}, /* 0x91d6 */
            {8'h00}, /* 0x91d5 */
            {8'h00}, /* 0x91d4 */
            {8'h00}, /* 0x91d3 */
            {8'h00}, /* 0x91d2 */
            {8'h00}, /* 0x91d1 */
            {8'h00}, /* 0x91d0 */
            {8'h00}, /* 0x91cf */
            {8'h00}, /* 0x91ce */
            {8'h00}, /* 0x91cd */
            {8'h00}, /* 0x91cc */
            {8'h00}, /* 0x91cb */
            {8'h00}, /* 0x91ca */
            {8'h00}, /* 0x91c9 */
            {8'h00}, /* 0x91c8 */
            {8'h00}, /* 0x91c7 */
            {8'h00}, /* 0x91c6 */
            {8'h00}, /* 0x91c5 */
            {8'h00}, /* 0x91c4 */
            {8'h00}, /* 0x91c3 */
            {8'h00}, /* 0x91c2 */
            {8'h00}, /* 0x91c1 */
            {8'h00}, /* 0x91c0 */
            {8'h00}, /* 0x91bf */
            {8'h00}, /* 0x91be */
            {8'h00}, /* 0x91bd */
            {8'h00}, /* 0x91bc */
            {8'h00}, /* 0x91bb */
            {8'h00}, /* 0x91ba */
            {8'h00}, /* 0x91b9 */
            {8'h00}, /* 0x91b8 */
            {8'h00}, /* 0x91b7 */
            {8'h00}, /* 0x91b6 */
            {8'h00}, /* 0x91b5 */
            {8'h00}, /* 0x91b4 */
            {8'h00}, /* 0x91b3 */
            {8'h00}, /* 0x91b2 */
            {8'h00}, /* 0x91b1 */
            {8'h00}, /* 0x91b0 */
            {8'h00}, /* 0x91af */
            {8'h00}, /* 0x91ae */
            {8'h00}, /* 0x91ad */
            {8'h00}, /* 0x91ac */
            {8'h00}, /* 0x91ab */
            {8'h00}, /* 0x91aa */
            {8'h00}, /* 0x91a9 */
            {8'h00}, /* 0x91a8 */
            {8'h00}, /* 0x91a7 */
            {8'h00}, /* 0x91a6 */
            {8'h00}, /* 0x91a5 */
            {8'h00}, /* 0x91a4 */
            {8'h00}, /* 0x91a3 */
            {8'h00}, /* 0x91a2 */
            {8'h00}, /* 0x91a1 */
            {8'h00}, /* 0x91a0 */
            {8'h00}, /* 0x919f */
            {8'h00}, /* 0x919e */
            {8'h00}, /* 0x919d */
            {8'h00}, /* 0x919c */
            {8'h00}, /* 0x919b */
            {8'h00}, /* 0x919a */
            {8'h00}, /* 0x9199 */
            {8'h00}, /* 0x9198 */
            {8'h00}, /* 0x9197 */
            {8'h00}, /* 0x9196 */
            {8'h00}, /* 0x9195 */
            {8'h00}, /* 0x9194 */
            {8'h00}, /* 0x9193 */
            {8'h00}, /* 0x9192 */
            {8'h00}, /* 0x9191 */
            {8'h00}, /* 0x9190 */
            {8'h00}, /* 0x918f */
            {8'h00}, /* 0x918e */
            {8'h00}, /* 0x918d */
            {8'h00}, /* 0x918c */
            {8'h00}, /* 0x918b */
            {8'h00}, /* 0x918a */
            {8'h00}, /* 0x9189 */
            {8'h00}, /* 0x9188 */
            {8'h00}, /* 0x9187 */
            {8'h00}, /* 0x9186 */
            {8'h00}, /* 0x9185 */
            {8'h00}, /* 0x9184 */
            {8'h00}, /* 0x9183 */
            {8'h00}, /* 0x9182 */
            {8'h00}, /* 0x9181 */
            {8'h00}, /* 0x9180 */
            {8'h00}, /* 0x917f */
            {8'h00}, /* 0x917e */
            {8'h00}, /* 0x917d */
            {8'h00}, /* 0x917c */
            {8'h00}, /* 0x917b */
            {8'h00}, /* 0x917a */
            {8'h00}, /* 0x9179 */
            {8'h00}, /* 0x9178 */
            {8'h00}, /* 0x9177 */
            {8'h00}, /* 0x9176 */
            {8'h00}, /* 0x9175 */
            {8'h00}, /* 0x9174 */
            {8'h00}, /* 0x9173 */
            {8'h00}, /* 0x9172 */
            {8'h00}, /* 0x9171 */
            {8'h00}, /* 0x9170 */
            {8'h00}, /* 0x916f */
            {8'h00}, /* 0x916e */
            {8'h00}, /* 0x916d */
            {8'h00}, /* 0x916c */
            {8'h00}, /* 0x916b */
            {8'h00}, /* 0x916a */
            {8'h00}, /* 0x9169 */
            {8'h00}, /* 0x9168 */
            {8'h00}, /* 0x9167 */
            {8'h00}, /* 0x9166 */
            {8'h00}, /* 0x9165 */
            {8'h00}, /* 0x9164 */
            {8'h00}, /* 0x9163 */
            {8'h00}, /* 0x9162 */
            {8'h00}, /* 0x9161 */
            {8'h00}, /* 0x9160 */
            {8'h00}, /* 0x915f */
            {8'h00}, /* 0x915e */
            {8'h00}, /* 0x915d */
            {8'h00}, /* 0x915c */
            {8'h00}, /* 0x915b */
            {8'h00}, /* 0x915a */
            {8'h00}, /* 0x9159 */
            {8'h00}, /* 0x9158 */
            {8'h00}, /* 0x9157 */
            {8'h00}, /* 0x9156 */
            {8'h00}, /* 0x9155 */
            {8'h00}, /* 0x9154 */
            {8'h00}, /* 0x9153 */
            {8'h00}, /* 0x9152 */
            {8'h00}, /* 0x9151 */
            {8'h00}, /* 0x9150 */
            {8'h00}, /* 0x914f */
            {8'h00}, /* 0x914e */
            {8'h00}, /* 0x914d */
            {8'h00}, /* 0x914c */
            {8'h00}, /* 0x914b */
            {8'h00}, /* 0x914a */
            {8'h00}, /* 0x9149 */
            {8'h00}, /* 0x9148 */
            {8'h00}, /* 0x9147 */
            {8'h00}, /* 0x9146 */
            {8'h00}, /* 0x9145 */
            {8'h00}, /* 0x9144 */
            {8'h00}, /* 0x9143 */
            {8'h00}, /* 0x9142 */
            {8'h00}, /* 0x9141 */
            {8'h00}, /* 0x9140 */
            {8'h00}, /* 0x913f */
            {8'h00}, /* 0x913e */
            {8'h00}, /* 0x913d */
            {8'h00}, /* 0x913c */
            {8'h00}, /* 0x913b */
            {8'h00}, /* 0x913a */
            {8'h00}, /* 0x9139 */
            {8'h00}, /* 0x9138 */
            {8'h00}, /* 0x9137 */
            {8'h00}, /* 0x9136 */
            {8'h00}, /* 0x9135 */
            {8'h00}, /* 0x9134 */
            {8'h00}, /* 0x9133 */
            {8'h00}, /* 0x9132 */
            {8'h00}, /* 0x9131 */
            {8'h00}, /* 0x9130 */
            {8'h00}, /* 0x912f */
            {8'h00}, /* 0x912e */
            {8'h00}, /* 0x912d */
            {8'h00}, /* 0x912c */
            {8'h00}, /* 0x912b */
            {8'h00}, /* 0x912a */
            {8'h00}, /* 0x9129 */
            {8'h00}, /* 0x9128 */
            {8'h00}, /* 0x9127 */
            {8'h00}, /* 0x9126 */
            {8'h00}, /* 0x9125 */
            {8'h00}, /* 0x9124 */
            {8'h00}, /* 0x9123 */
            {8'h00}, /* 0x9122 */
            {8'h00}, /* 0x9121 */
            {8'h00}, /* 0x9120 */
            {8'h00}, /* 0x911f */
            {8'h00}, /* 0x911e */
            {8'h00}, /* 0x911d */
            {8'h00}, /* 0x911c */
            {8'h00}, /* 0x911b */
            {8'h00}, /* 0x911a */
            {8'h00}, /* 0x9119 */
            {8'h00}, /* 0x9118 */
            {8'h00}, /* 0x9117 */
            {8'h00}, /* 0x9116 */
            {8'h00}, /* 0x9115 */
            {8'h00}, /* 0x9114 */
            {8'h00}, /* 0x9113 */
            {8'h00}, /* 0x9112 */
            {8'h00}, /* 0x9111 */
            {8'h00}, /* 0x9110 */
            {8'h00}, /* 0x910f */
            {8'h00}, /* 0x910e */
            {8'h00}, /* 0x910d */
            {8'h00}, /* 0x910c */
            {8'h00}, /* 0x910b */
            {8'h00}, /* 0x910a */
            {8'h00}, /* 0x9109 */
            {8'h00}, /* 0x9108 */
            {8'h00}, /* 0x9107 */
            {8'h00}, /* 0x9106 */
            {8'h00}, /* 0x9105 */
            {8'h00}, /* 0x9104 */
            {8'h00}, /* 0x9103 */
            {8'h00}, /* 0x9102 */
            {8'h00}, /* 0x9101 */
            {8'h00}, /* 0x9100 */
            {8'h00}, /* 0x90ff */
            {8'h00}, /* 0x90fe */
            {8'h00}, /* 0x90fd */
            {8'h00}, /* 0x90fc */
            {8'h00}, /* 0x90fb */
            {8'h00}, /* 0x90fa */
            {8'h00}, /* 0x90f9 */
            {8'h00}, /* 0x90f8 */
            {8'h00}, /* 0x90f7 */
            {8'h00}, /* 0x90f6 */
            {8'h00}, /* 0x90f5 */
            {8'h00}, /* 0x90f4 */
            {8'h00}, /* 0x90f3 */
            {8'h00}, /* 0x90f2 */
            {8'h00}, /* 0x90f1 */
            {8'h00}, /* 0x90f0 */
            {8'h00}, /* 0x90ef */
            {8'h00}, /* 0x90ee */
            {8'h00}, /* 0x90ed */
            {8'h00}, /* 0x90ec */
            {8'h00}, /* 0x90eb */
            {8'h00}, /* 0x90ea */
            {8'h00}, /* 0x90e9 */
            {8'h00}, /* 0x90e8 */
            {8'h00}, /* 0x90e7 */
            {8'h00}, /* 0x90e6 */
            {8'h00}, /* 0x90e5 */
            {8'h00}, /* 0x90e4 */
            {8'h00}, /* 0x90e3 */
            {8'h00}, /* 0x90e2 */
            {8'h00}, /* 0x90e1 */
            {8'h00}, /* 0x90e0 */
            {8'h00}, /* 0x90df */
            {8'h00}, /* 0x90de */
            {8'h00}, /* 0x90dd */
            {8'h00}, /* 0x90dc */
            {8'h00}, /* 0x90db */
            {8'h00}, /* 0x90da */
            {8'h00}, /* 0x90d9 */
            {8'h00}, /* 0x90d8 */
            {8'h00}, /* 0x90d7 */
            {8'h00}, /* 0x90d6 */
            {8'h00}, /* 0x90d5 */
            {8'h00}, /* 0x90d4 */
            {8'h00}, /* 0x90d3 */
            {8'h00}, /* 0x90d2 */
            {8'h00}, /* 0x90d1 */
            {8'h00}, /* 0x90d0 */
            {8'h00}, /* 0x90cf */
            {8'h00}, /* 0x90ce */
            {8'h00}, /* 0x90cd */
            {8'h00}, /* 0x90cc */
            {8'h00}, /* 0x90cb */
            {8'h00}, /* 0x90ca */
            {8'h00}, /* 0x90c9 */
            {8'h00}, /* 0x90c8 */
            {8'h00}, /* 0x90c7 */
            {8'h00}, /* 0x90c6 */
            {8'h00}, /* 0x90c5 */
            {8'h00}, /* 0x90c4 */
            {8'h00}, /* 0x90c3 */
            {8'h00}, /* 0x90c2 */
            {8'h00}, /* 0x90c1 */
            {8'h00}, /* 0x90c0 */
            {8'h00}, /* 0x90bf */
            {8'h00}, /* 0x90be */
            {8'h00}, /* 0x90bd */
            {8'h00}, /* 0x90bc */
            {8'h00}, /* 0x90bb */
            {8'h00}, /* 0x90ba */
            {8'h00}, /* 0x90b9 */
            {8'h00}, /* 0x90b8 */
            {8'h00}, /* 0x90b7 */
            {8'h00}, /* 0x90b6 */
            {8'h00}, /* 0x90b5 */
            {8'h00}, /* 0x90b4 */
            {8'h00}, /* 0x90b3 */
            {8'h00}, /* 0x90b2 */
            {8'h00}, /* 0x90b1 */
            {8'h00}, /* 0x90b0 */
            {8'h00}, /* 0x90af */
            {8'h00}, /* 0x90ae */
            {8'h00}, /* 0x90ad */
            {8'h00}, /* 0x90ac */
            {8'h00}, /* 0x90ab */
            {8'h00}, /* 0x90aa */
            {8'h00}, /* 0x90a9 */
            {8'h00}, /* 0x90a8 */
            {8'h00}, /* 0x90a7 */
            {8'h00}, /* 0x90a6 */
            {8'h00}, /* 0x90a5 */
            {8'h00}, /* 0x90a4 */
            {8'h00}, /* 0x90a3 */
            {8'h00}, /* 0x90a2 */
            {8'h00}, /* 0x90a1 */
            {8'h00}, /* 0x90a0 */
            {8'h00}, /* 0x909f */
            {8'h00}, /* 0x909e */
            {8'h00}, /* 0x909d */
            {8'h00}, /* 0x909c */
            {8'h00}, /* 0x909b */
            {8'h00}, /* 0x909a */
            {8'h00}, /* 0x9099 */
            {8'h00}, /* 0x9098 */
            {8'h00}, /* 0x9097 */
            {8'h00}, /* 0x9096 */
            {8'h00}, /* 0x9095 */
            {8'h00}, /* 0x9094 */
            {8'h00}, /* 0x9093 */
            {8'h00}, /* 0x9092 */
            {8'h00}, /* 0x9091 */
            {8'h00}, /* 0x9090 */
            {8'h00}, /* 0x908f */
            {8'h00}, /* 0x908e */
            {8'h00}, /* 0x908d */
            {8'h00}, /* 0x908c */
            {8'h00}, /* 0x908b */
            {8'h00}, /* 0x908a */
            {8'h00}, /* 0x9089 */
            {8'h00}, /* 0x9088 */
            {8'h00}, /* 0x9087 */
            {8'h00}, /* 0x9086 */
            {8'h00}, /* 0x9085 */
            {8'h00}, /* 0x9084 */
            {8'h00}, /* 0x9083 */
            {8'h00}, /* 0x9082 */
            {8'h00}, /* 0x9081 */
            {8'h00}, /* 0x9080 */
            {8'h00}, /* 0x907f */
            {8'h00}, /* 0x907e */
            {8'h00}, /* 0x907d */
            {8'h00}, /* 0x907c */
            {8'h00}, /* 0x907b */
            {8'h00}, /* 0x907a */
            {8'h00}, /* 0x9079 */
            {8'h00}, /* 0x9078 */
            {8'h00}, /* 0x9077 */
            {8'h00}, /* 0x9076 */
            {8'h00}, /* 0x9075 */
            {8'h00}, /* 0x9074 */
            {8'h00}, /* 0x9073 */
            {8'h00}, /* 0x9072 */
            {8'h00}, /* 0x9071 */
            {8'h00}, /* 0x9070 */
            {8'h00}, /* 0x906f */
            {8'h00}, /* 0x906e */
            {8'h00}, /* 0x906d */
            {8'h00}, /* 0x906c */
            {8'h00}, /* 0x906b */
            {8'h00}, /* 0x906a */
            {8'h00}, /* 0x9069 */
            {8'h00}, /* 0x9068 */
            {8'h00}, /* 0x9067 */
            {8'h00}, /* 0x9066 */
            {8'h00}, /* 0x9065 */
            {8'h00}, /* 0x9064 */
            {8'h00}, /* 0x9063 */
            {8'h00}, /* 0x9062 */
            {8'h00}, /* 0x9061 */
            {8'h00}, /* 0x9060 */
            {8'h00}, /* 0x905f */
            {8'h00}, /* 0x905e */
            {8'h00}, /* 0x905d */
            {8'h00}, /* 0x905c */
            {8'h00}, /* 0x905b */
            {8'h00}, /* 0x905a */
            {8'h00}, /* 0x9059 */
            {8'h00}, /* 0x9058 */
            {8'h00}, /* 0x9057 */
            {8'h00}, /* 0x9056 */
            {8'h00}, /* 0x9055 */
            {8'h00}, /* 0x9054 */
            {8'h00}, /* 0x9053 */
            {8'h00}, /* 0x9052 */
            {8'h00}, /* 0x9051 */
            {8'h00}, /* 0x9050 */
            {8'h00}, /* 0x904f */
            {8'h00}, /* 0x904e */
            {8'h00}, /* 0x904d */
            {8'h00}, /* 0x904c */
            {8'h00}, /* 0x904b */
            {8'h00}, /* 0x904a */
            {8'h00}, /* 0x9049 */
            {8'h00}, /* 0x9048 */
            {8'h00}, /* 0x9047 */
            {8'h00}, /* 0x9046 */
            {8'h00}, /* 0x9045 */
            {8'h00}, /* 0x9044 */
            {8'h00}, /* 0x9043 */
            {8'h00}, /* 0x9042 */
            {8'h00}, /* 0x9041 */
            {8'h00}, /* 0x9040 */
            {8'h00}, /* 0x903f */
            {8'h00}, /* 0x903e */
            {8'h00}, /* 0x903d */
            {8'h00}, /* 0x903c */
            {8'h00}, /* 0x903b */
            {8'h00}, /* 0x903a */
            {8'h00}, /* 0x9039 */
            {8'h00}, /* 0x9038 */
            {8'h00}, /* 0x9037 */
            {8'h00}, /* 0x9036 */
            {8'h00}, /* 0x9035 */
            {8'h00}, /* 0x9034 */
            {8'h00}, /* 0x9033 */
            {8'h00}, /* 0x9032 */
            {8'h00}, /* 0x9031 */
            {8'h00}, /* 0x9030 */
            {8'h00}, /* 0x902f */
            {8'h00}, /* 0x902e */
            {8'h00}, /* 0x902d */
            {8'h00}, /* 0x902c */
            {8'h00}, /* 0x902b */
            {8'h00}, /* 0x902a */
            {8'h00}, /* 0x9029 */
            {8'h00}, /* 0x9028 */
            {8'h00}, /* 0x9027 */
            {8'h00}, /* 0x9026 */
            {8'h00}, /* 0x9025 */
            {8'h00}, /* 0x9024 */
            {8'h00}, /* 0x9023 */
            {8'h00}, /* 0x9022 */
            {8'h00}, /* 0x9021 */
            {8'h00}, /* 0x9020 */
            {8'h00}, /* 0x901f */
            {8'h00}, /* 0x901e */
            {8'h00}, /* 0x901d */
            {8'h00}, /* 0x901c */
            {8'h00}, /* 0x901b */
            {8'h00}, /* 0x901a */
            {8'h00}, /* 0x9019 */
            {8'h00}, /* 0x9018 */
            {8'h00}, /* 0x9017 */
            {8'h00}, /* 0x9016 */
            {8'h00}, /* 0x9015 */
            {8'h00}, /* 0x9014 */
            {8'h00}, /* 0x9013 */
            {8'h00}, /* 0x9012 */
            {8'h00}, /* 0x9011 */
            {8'h00}, /* 0x9010 */
            {8'h00}, /* 0x900f */
            {8'h00}, /* 0x900e */
            {8'h00}, /* 0x900d */
            {8'h00}, /* 0x900c */
            {8'h00}, /* 0x900b */
            {8'h00}, /* 0x900a */
            {8'h00}, /* 0x9009 */
            {8'h00}, /* 0x9008 */
            {8'h00}, /* 0x9007 */
            {8'h00}, /* 0x9006 */
            {8'h00}, /* 0x9005 */
            {8'h00}, /* 0x9004 */
            {8'h00}, /* 0x9003 */
            {8'h00}, /* 0x9002 */
            {8'h00}, /* 0x9001 */
            {8'h00}, /* 0x9000 */
            {8'h00}, /* 0x8fff */
            {8'h00}, /* 0x8ffe */
            {8'h00}, /* 0x8ffd */
            {8'h00}, /* 0x8ffc */
            {8'h00}, /* 0x8ffb */
            {8'h00}, /* 0x8ffa */
            {8'h00}, /* 0x8ff9 */
            {8'h00}, /* 0x8ff8 */
            {8'h00}, /* 0x8ff7 */
            {8'h00}, /* 0x8ff6 */
            {8'h00}, /* 0x8ff5 */
            {8'h00}, /* 0x8ff4 */
            {8'h00}, /* 0x8ff3 */
            {8'h00}, /* 0x8ff2 */
            {8'h00}, /* 0x8ff1 */
            {8'h00}, /* 0x8ff0 */
            {8'h00}, /* 0x8fef */
            {8'h00}, /* 0x8fee */
            {8'h00}, /* 0x8fed */
            {8'h00}, /* 0x8fec */
            {8'h00}, /* 0x8feb */
            {8'h00}, /* 0x8fea */
            {8'h00}, /* 0x8fe9 */
            {8'h00}, /* 0x8fe8 */
            {8'h00}, /* 0x8fe7 */
            {8'h00}, /* 0x8fe6 */
            {8'h00}, /* 0x8fe5 */
            {8'h00}, /* 0x8fe4 */
            {8'h00}, /* 0x8fe3 */
            {8'h00}, /* 0x8fe2 */
            {8'h00}, /* 0x8fe1 */
            {8'h00}, /* 0x8fe0 */
            {8'h00}, /* 0x8fdf */
            {8'h00}, /* 0x8fde */
            {8'h00}, /* 0x8fdd */
            {8'h00}, /* 0x8fdc */
            {8'h00}, /* 0x8fdb */
            {8'h00}, /* 0x8fda */
            {8'h00}, /* 0x8fd9 */
            {8'h00}, /* 0x8fd8 */
            {8'h00}, /* 0x8fd7 */
            {8'h00}, /* 0x8fd6 */
            {8'h00}, /* 0x8fd5 */
            {8'h00}, /* 0x8fd4 */
            {8'h00}, /* 0x8fd3 */
            {8'h00}, /* 0x8fd2 */
            {8'h00}, /* 0x8fd1 */
            {8'h00}, /* 0x8fd0 */
            {8'h00}, /* 0x8fcf */
            {8'h00}, /* 0x8fce */
            {8'h00}, /* 0x8fcd */
            {8'h00}, /* 0x8fcc */
            {8'h00}, /* 0x8fcb */
            {8'h00}, /* 0x8fca */
            {8'h00}, /* 0x8fc9 */
            {8'h00}, /* 0x8fc8 */
            {8'h00}, /* 0x8fc7 */
            {8'h00}, /* 0x8fc6 */
            {8'h00}, /* 0x8fc5 */
            {8'h00}, /* 0x8fc4 */
            {8'h00}, /* 0x8fc3 */
            {8'h00}, /* 0x8fc2 */
            {8'h00}, /* 0x8fc1 */
            {8'h00}, /* 0x8fc0 */
            {8'h00}, /* 0x8fbf */
            {8'h00}, /* 0x8fbe */
            {8'h00}, /* 0x8fbd */
            {8'h00}, /* 0x8fbc */
            {8'h00}, /* 0x8fbb */
            {8'h00}, /* 0x8fba */
            {8'h00}, /* 0x8fb9 */
            {8'h00}, /* 0x8fb8 */
            {8'h00}, /* 0x8fb7 */
            {8'h00}, /* 0x8fb6 */
            {8'h00}, /* 0x8fb5 */
            {8'h00}, /* 0x8fb4 */
            {8'h00}, /* 0x8fb3 */
            {8'h00}, /* 0x8fb2 */
            {8'h00}, /* 0x8fb1 */
            {8'h00}, /* 0x8fb0 */
            {8'h00}, /* 0x8faf */
            {8'h00}, /* 0x8fae */
            {8'h00}, /* 0x8fad */
            {8'h00}, /* 0x8fac */
            {8'h00}, /* 0x8fab */
            {8'h00}, /* 0x8faa */
            {8'h00}, /* 0x8fa9 */
            {8'h00}, /* 0x8fa8 */
            {8'h00}, /* 0x8fa7 */
            {8'h00}, /* 0x8fa6 */
            {8'h00}, /* 0x8fa5 */
            {8'h00}, /* 0x8fa4 */
            {8'h00}, /* 0x8fa3 */
            {8'h00}, /* 0x8fa2 */
            {8'h00}, /* 0x8fa1 */
            {8'h00}, /* 0x8fa0 */
            {8'h00}, /* 0x8f9f */
            {8'h00}, /* 0x8f9e */
            {8'h00}, /* 0x8f9d */
            {8'h00}, /* 0x8f9c */
            {8'h00}, /* 0x8f9b */
            {8'h00}, /* 0x8f9a */
            {8'h00}, /* 0x8f99 */
            {8'h00}, /* 0x8f98 */
            {8'h00}, /* 0x8f97 */
            {8'h00}, /* 0x8f96 */
            {8'h00}, /* 0x8f95 */
            {8'h00}, /* 0x8f94 */
            {8'h00}, /* 0x8f93 */
            {8'h00}, /* 0x8f92 */
            {8'h00}, /* 0x8f91 */
            {8'h00}, /* 0x8f90 */
            {8'h00}, /* 0x8f8f */
            {8'h00}, /* 0x8f8e */
            {8'h00}, /* 0x8f8d */
            {8'h00}, /* 0x8f8c */
            {8'h00}, /* 0x8f8b */
            {8'h00}, /* 0x8f8a */
            {8'h00}, /* 0x8f89 */
            {8'h00}, /* 0x8f88 */
            {8'h00}, /* 0x8f87 */
            {8'h00}, /* 0x8f86 */
            {8'h00}, /* 0x8f85 */
            {8'h00}, /* 0x8f84 */
            {8'h00}, /* 0x8f83 */
            {8'h00}, /* 0x8f82 */
            {8'h00}, /* 0x8f81 */
            {8'h00}, /* 0x8f80 */
            {8'h00}, /* 0x8f7f */
            {8'h00}, /* 0x8f7e */
            {8'h00}, /* 0x8f7d */
            {8'h00}, /* 0x8f7c */
            {8'h00}, /* 0x8f7b */
            {8'h00}, /* 0x8f7a */
            {8'h00}, /* 0x8f79 */
            {8'h00}, /* 0x8f78 */
            {8'h00}, /* 0x8f77 */
            {8'h00}, /* 0x8f76 */
            {8'h00}, /* 0x8f75 */
            {8'h00}, /* 0x8f74 */
            {8'h00}, /* 0x8f73 */
            {8'h00}, /* 0x8f72 */
            {8'h00}, /* 0x8f71 */
            {8'h00}, /* 0x8f70 */
            {8'h00}, /* 0x8f6f */
            {8'h00}, /* 0x8f6e */
            {8'h00}, /* 0x8f6d */
            {8'h00}, /* 0x8f6c */
            {8'h00}, /* 0x8f6b */
            {8'h00}, /* 0x8f6a */
            {8'h00}, /* 0x8f69 */
            {8'h00}, /* 0x8f68 */
            {8'h00}, /* 0x8f67 */
            {8'h00}, /* 0x8f66 */
            {8'h00}, /* 0x8f65 */
            {8'h00}, /* 0x8f64 */
            {8'h00}, /* 0x8f63 */
            {8'h00}, /* 0x8f62 */
            {8'h00}, /* 0x8f61 */
            {8'h00}, /* 0x8f60 */
            {8'h00}, /* 0x8f5f */
            {8'h00}, /* 0x8f5e */
            {8'h00}, /* 0x8f5d */
            {8'h00}, /* 0x8f5c */
            {8'h00}, /* 0x8f5b */
            {8'h00}, /* 0x8f5a */
            {8'h00}, /* 0x8f59 */
            {8'h00}, /* 0x8f58 */
            {8'h00}, /* 0x8f57 */
            {8'h00}, /* 0x8f56 */
            {8'h00}, /* 0x8f55 */
            {8'h00}, /* 0x8f54 */
            {8'h00}, /* 0x8f53 */
            {8'h00}, /* 0x8f52 */
            {8'h00}, /* 0x8f51 */
            {8'h00}, /* 0x8f50 */
            {8'h00}, /* 0x8f4f */
            {8'h00}, /* 0x8f4e */
            {8'h00}, /* 0x8f4d */
            {8'h00}, /* 0x8f4c */
            {8'h00}, /* 0x8f4b */
            {8'h00}, /* 0x8f4a */
            {8'h00}, /* 0x8f49 */
            {8'h00}, /* 0x8f48 */
            {8'h00}, /* 0x8f47 */
            {8'h00}, /* 0x8f46 */
            {8'h00}, /* 0x8f45 */
            {8'h00}, /* 0x8f44 */
            {8'h00}, /* 0x8f43 */
            {8'h00}, /* 0x8f42 */
            {8'h00}, /* 0x8f41 */
            {8'h00}, /* 0x8f40 */
            {8'h00}, /* 0x8f3f */
            {8'h00}, /* 0x8f3e */
            {8'h00}, /* 0x8f3d */
            {8'h00}, /* 0x8f3c */
            {8'h00}, /* 0x8f3b */
            {8'h00}, /* 0x8f3a */
            {8'h00}, /* 0x8f39 */
            {8'h00}, /* 0x8f38 */
            {8'h00}, /* 0x8f37 */
            {8'h00}, /* 0x8f36 */
            {8'h00}, /* 0x8f35 */
            {8'h00}, /* 0x8f34 */
            {8'h00}, /* 0x8f33 */
            {8'h00}, /* 0x8f32 */
            {8'h00}, /* 0x8f31 */
            {8'h00}, /* 0x8f30 */
            {8'h00}, /* 0x8f2f */
            {8'h00}, /* 0x8f2e */
            {8'h00}, /* 0x8f2d */
            {8'h00}, /* 0x8f2c */
            {8'h00}, /* 0x8f2b */
            {8'h00}, /* 0x8f2a */
            {8'h00}, /* 0x8f29 */
            {8'h00}, /* 0x8f28 */
            {8'h00}, /* 0x8f27 */
            {8'h00}, /* 0x8f26 */
            {8'h00}, /* 0x8f25 */
            {8'h00}, /* 0x8f24 */
            {8'h00}, /* 0x8f23 */
            {8'h00}, /* 0x8f22 */
            {8'h00}, /* 0x8f21 */
            {8'h00}, /* 0x8f20 */
            {8'h00}, /* 0x8f1f */
            {8'h00}, /* 0x8f1e */
            {8'h00}, /* 0x8f1d */
            {8'h00}, /* 0x8f1c */
            {8'h00}, /* 0x8f1b */
            {8'h00}, /* 0x8f1a */
            {8'h00}, /* 0x8f19 */
            {8'h00}, /* 0x8f18 */
            {8'h00}, /* 0x8f17 */
            {8'h00}, /* 0x8f16 */
            {8'h00}, /* 0x8f15 */
            {8'h00}, /* 0x8f14 */
            {8'h00}, /* 0x8f13 */
            {8'h00}, /* 0x8f12 */
            {8'h00}, /* 0x8f11 */
            {8'h00}, /* 0x8f10 */
            {8'h00}, /* 0x8f0f */
            {8'h00}, /* 0x8f0e */
            {8'h00}, /* 0x8f0d */
            {8'h00}, /* 0x8f0c */
            {8'h00}, /* 0x8f0b */
            {8'h00}, /* 0x8f0a */
            {8'h00}, /* 0x8f09 */
            {8'h00}, /* 0x8f08 */
            {8'h00}, /* 0x8f07 */
            {8'h00}, /* 0x8f06 */
            {8'h00}, /* 0x8f05 */
            {8'h00}, /* 0x8f04 */
            {8'h00}, /* 0x8f03 */
            {8'h00}, /* 0x8f02 */
            {8'h00}, /* 0x8f01 */
            {8'h00}, /* 0x8f00 */
            {8'h00}, /* 0x8eff */
            {8'h00}, /* 0x8efe */
            {8'h00}, /* 0x8efd */
            {8'h00}, /* 0x8efc */
            {8'h00}, /* 0x8efb */
            {8'h00}, /* 0x8efa */
            {8'h00}, /* 0x8ef9 */
            {8'h00}, /* 0x8ef8 */
            {8'h00}, /* 0x8ef7 */
            {8'h00}, /* 0x8ef6 */
            {8'h00}, /* 0x8ef5 */
            {8'h00}, /* 0x8ef4 */
            {8'h00}, /* 0x8ef3 */
            {8'h00}, /* 0x8ef2 */
            {8'h00}, /* 0x8ef1 */
            {8'h00}, /* 0x8ef0 */
            {8'h00}, /* 0x8eef */
            {8'h00}, /* 0x8eee */
            {8'h00}, /* 0x8eed */
            {8'h00}, /* 0x8eec */
            {8'h00}, /* 0x8eeb */
            {8'h00}, /* 0x8eea */
            {8'h00}, /* 0x8ee9 */
            {8'h00}, /* 0x8ee8 */
            {8'h00}, /* 0x8ee7 */
            {8'h00}, /* 0x8ee6 */
            {8'h00}, /* 0x8ee5 */
            {8'h00}, /* 0x8ee4 */
            {8'h00}, /* 0x8ee3 */
            {8'h00}, /* 0x8ee2 */
            {8'h00}, /* 0x8ee1 */
            {8'h00}, /* 0x8ee0 */
            {8'h00}, /* 0x8edf */
            {8'h00}, /* 0x8ede */
            {8'h00}, /* 0x8edd */
            {8'h00}, /* 0x8edc */
            {8'h00}, /* 0x8edb */
            {8'h00}, /* 0x8eda */
            {8'h00}, /* 0x8ed9 */
            {8'h00}, /* 0x8ed8 */
            {8'h00}, /* 0x8ed7 */
            {8'h00}, /* 0x8ed6 */
            {8'h00}, /* 0x8ed5 */
            {8'h00}, /* 0x8ed4 */
            {8'h00}, /* 0x8ed3 */
            {8'h00}, /* 0x8ed2 */
            {8'h00}, /* 0x8ed1 */
            {8'h00}, /* 0x8ed0 */
            {8'h00}, /* 0x8ecf */
            {8'h00}, /* 0x8ece */
            {8'h00}, /* 0x8ecd */
            {8'h00}, /* 0x8ecc */
            {8'h00}, /* 0x8ecb */
            {8'h00}, /* 0x8eca */
            {8'h00}, /* 0x8ec9 */
            {8'h00}, /* 0x8ec8 */
            {8'h00}, /* 0x8ec7 */
            {8'h00}, /* 0x8ec6 */
            {8'h00}, /* 0x8ec5 */
            {8'h00}, /* 0x8ec4 */
            {8'h00}, /* 0x8ec3 */
            {8'h00}, /* 0x8ec2 */
            {8'h00}, /* 0x8ec1 */
            {8'h00}, /* 0x8ec0 */
            {8'h00}, /* 0x8ebf */
            {8'h00}, /* 0x8ebe */
            {8'h00}, /* 0x8ebd */
            {8'h00}, /* 0x8ebc */
            {8'h00}, /* 0x8ebb */
            {8'h00}, /* 0x8eba */
            {8'h00}, /* 0x8eb9 */
            {8'h00}, /* 0x8eb8 */
            {8'h00}, /* 0x8eb7 */
            {8'h00}, /* 0x8eb6 */
            {8'h00}, /* 0x8eb5 */
            {8'h00}, /* 0x8eb4 */
            {8'h00}, /* 0x8eb3 */
            {8'h00}, /* 0x8eb2 */
            {8'h00}, /* 0x8eb1 */
            {8'h00}, /* 0x8eb0 */
            {8'h00}, /* 0x8eaf */
            {8'h00}, /* 0x8eae */
            {8'h00}, /* 0x8ead */
            {8'h00}, /* 0x8eac */
            {8'h00}, /* 0x8eab */
            {8'h00}, /* 0x8eaa */
            {8'h00}, /* 0x8ea9 */
            {8'h00}, /* 0x8ea8 */
            {8'h00}, /* 0x8ea7 */
            {8'h00}, /* 0x8ea6 */
            {8'h00}, /* 0x8ea5 */
            {8'h00}, /* 0x8ea4 */
            {8'h00}, /* 0x8ea3 */
            {8'h00}, /* 0x8ea2 */
            {8'h00}, /* 0x8ea1 */
            {8'h00}, /* 0x8ea0 */
            {8'h00}, /* 0x8e9f */
            {8'h00}, /* 0x8e9e */
            {8'h00}, /* 0x8e9d */
            {8'h00}, /* 0x8e9c */
            {8'h00}, /* 0x8e9b */
            {8'h00}, /* 0x8e9a */
            {8'h00}, /* 0x8e99 */
            {8'h00}, /* 0x8e98 */
            {8'h00}, /* 0x8e97 */
            {8'h00}, /* 0x8e96 */
            {8'h00}, /* 0x8e95 */
            {8'h00}, /* 0x8e94 */
            {8'h00}, /* 0x8e93 */
            {8'h00}, /* 0x8e92 */
            {8'h00}, /* 0x8e91 */
            {8'h00}, /* 0x8e90 */
            {8'h00}, /* 0x8e8f */
            {8'h00}, /* 0x8e8e */
            {8'h00}, /* 0x8e8d */
            {8'h00}, /* 0x8e8c */
            {8'h00}, /* 0x8e8b */
            {8'h00}, /* 0x8e8a */
            {8'h00}, /* 0x8e89 */
            {8'h00}, /* 0x8e88 */
            {8'h00}, /* 0x8e87 */
            {8'h00}, /* 0x8e86 */
            {8'h00}, /* 0x8e85 */
            {8'h00}, /* 0x8e84 */
            {8'h00}, /* 0x8e83 */
            {8'h00}, /* 0x8e82 */
            {8'h00}, /* 0x8e81 */
            {8'h00}, /* 0x8e80 */
            {8'h00}, /* 0x8e7f */
            {8'h00}, /* 0x8e7e */
            {8'h00}, /* 0x8e7d */
            {8'h00}, /* 0x8e7c */
            {8'h00}, /* 0x8e7b */
            {8'h00}, /* 0x8e7a */
            {8'h00}, /* 0x8e79 */
            {8'h00}, /* 0x8e78 */
            {8'h00}, /* 0x8e77 */
            {8'h00}, /* 0x8e76 */
            {8'h00}, /* 0x8e75 */
            {8'h00}, /* 0x8e74 */
            {8'h00}, /* 0x8e73 */
            {8'h00}, /* 0x8e72 */
            {8'h00}, /* 0x8e71 */
            {8'h00}, /* 0x8e70 */
            {8'h00}, /* 0x8e6f */
            {8'h00}, /* 0x8e6e */
            {8'h00}, /* 0x8e6d */
            {8'h00}, /* 0x8e6c */
            {8'h00}, /* 0x8e6b */
            {8'h00}, /* 0x8e6a */
            {8'h00}, /* 0x8e69 */
            {8'h00}, /* 0x8e68 */
            {8'h00}, /* 0x8e67 */
            {8'h00}, /* 0x8e66 */
            {8'h00}, /* 0x8e65 */
            {8'h00}, /* 0x8e64 */
            {8'h00}, /* 0x8e63 */
            {8'h00}, /* 0x8e62 */
            {8'h00}, /* 0x8e61 */
            {8'h00}, /* 0x8e60 */
            {8'h00}, /* 0x8e5f */
            {8'h00}, /* 0x8e5e */
            {8'h00}, /* 0x8e5d */
            {8'h00}, /* 0x8e5c */
            {8'h00}, /* 0x8e5b */
            {8'h00}, /* 0x8e5a */
            {8'h00}, /* 0x8e59 */
            {8'h00}, /* 0x8e58 */
            {8'h00}, /* 0x8e57 */
            {8'h00}, /* 0x8e56 */
            {8'h00}, /* 0x8e55 */
            {8'h00}, /* 0x8e54 */
            {8'h00}, /* 0x8e53 */
            {8'h00}, /* 0x8e52 */
            {8'h00}, /* 0x8e51 */
            {8'h00}, /* 0x8e50 */
            {8'h00}, /* 0x8e4f */
            {8'h00}, /* 0x8e4e */
            {8'h00}, /* 0x8e4d */
            {8'h00}, /* 0x8e4c */
            {8'h00}, /* 0x8e4b */
            {8'h00}, /* 0x8e4a */
            {8'h00}, /* 0x8e49 */
            {8'h00}, /* 0x8e48 */
            {8'h00}, /* 0x8e47 */
            {8'h00}, /* 0x8e46 */
            {8'h00}, /* 0x8e45 */
            {8'h00}, /* 0x8e44 */
            {8'h00}, /* 0x8e43 */
            {8'h00}, /* 0x8e42 */
            {8'h00}, /* 0x8e41 */
            {8'h00}, /* 0x8e40 */
            {8'h00}, /* 0x8e3f */
            {8'h00}, /* 0x8e3e */
            {8'h00}, /* 0x8e3d */
            {8'h00}, /* 0x8e3c */
            {8'h00}, /* 0x8e3b */
            {8'h00}, /* 0x8e3a */
            {8'h00}, /* 0x8e39 */
            {8'h00}, /* 0x8e38 */
            {8'h00}, /* 0x8e37 */
            {8'h00}, /* 0x8e36 */
            {8'h00}, /* 0x8e35 */
            {8'h00}, /* 0x8e34 */
            {8'h00}, /* 0x8e33 */
            {8'h00}, /* 0x8e32 */
            {8'h00}, /* 0x8e31 */
            {8'h00}, /* 0x8e30 */
            {8'h00}, /* 0x8e2f */
            {8'h00}, /* 0x8e2e */
            {8'h00}, /* 0x8e2d */
            {8'h00}, /* 0x8e2c */
            {8'h00}, /* 0x8e2b */
            {8'h00}, /* 0x8e2a */
            {8'h00}, /* 0x8e29 */
            {8'h00}, /* 0x8e28 */
            {8'h00}, /* 0x8e27 */
            {8'h00}, /* 0x8e26 */
            {8'h00}, /* 0x8e25 */
            {8'h00}, /* 0x8e24 */
            {8'h00}, /* 0x8e23 */
            {8'h00}, /* 0x8e22 */
            {8'h00}, /* 0x8e21 */
            {8'h00}, /* 0x8e20 */
            {8'h00}, /* 0x8e1f */
            {8'h00}, /* 0x8e1e */
            {8'h00}, /* 0x8e1d */
            {8'h00}, /* 0x8e1c */
            {8'h00}, /* 0x8e1b */
            {8'h00}, /* 0x8e1a */
            {8'h00}, /* 0x8e19 */
            {8'h00}, /* 0x8e18 */
            {8'h00}, /* 0x8e17 */
            {8'h00}, /* 0x8e16 */
            {8'h00}, /* 0x8e15 */
            {8'h00}, /* 0x8e14 */
            {8'h00}, /* 0x8e13 */
            {8'h00}, /* 0x8e12 */
            {8'h00}, /* 0x8e11 */
            {8'h00}, /* 0x8e10 */
            {8'h00}, /* 0x8e0f */
            {8'h00}, /* 0x8e0e */
            {8'h00}, /* 0x8e0d */
            {8'h00}, /* 0x8e0c */
            {8'h00}, /* 0x8e0b */
            {8'h00}, /* 0x8e0a */
            {8'h00}, /* 0x8e09 */
            {8'h00}, /* 0x8e08 */
            {8'h00}, /* 0x8e07 */
            {8'h00}, /* 0x8e06 */
            {8'h00}, /* 0x8e05 */
            {8'h00}, /* 0x8e04 */
            {8'h00}, /* 0x8e03 */
            {8'h00}, /* 0x8e02 */
            {8'h00}, /* 0x8e01 */
            {8'h00}, /* 0x8e00 */
            {8'h00}, /* 0x8dff */
            {8'h00}, /* 0x8dfe */
            {8'h00}, /* 0x8dfd */
            {8'h00}, /* 0x8dfc */
            {8'h00}, /* 0x8dfb */
            {8'h00}, /* 0x8dfa */
            {8'h00}, /* 0x8df9 */
            {8'h00}, /* 0x8df8 */
            {8'h00}, /* 0x8df7 */
            {8'h00}, /* 0x8df6 */
            {8'h00}, /* 0x8df5 */
            {8'h00}, /* 0x8df4 */
            {8'h00}, /* 0x8df3 */
            {8'h00}, /* 0x8df2 */
            {8'h00}, /* 0x8df1 */
            {8'h00}, /* 0x8df0 */
            {8'h00}, /* 0x8def */
            {8'h00}, /* 0x8dee */
            {8'h00}, /* 0x8ded */
            {8'h00}, /* 0x8dec */
            {8'h00}, /* 0x8deb */
            {8'h00}, /* 0x8dea */
            {8'h00}, /* 0x8de9 */
            {8'h00}, /* 0x8de8 */
            {8'h00}, /* 0x8de7 */
            {8'h00}, /* 0x8de6 */
            {8'h00}, /* 0x8de5 */
            {8'h00}, /* 0x8de4 */
            {8'h00}, /* 0x8de3 */
            {8'h00}, /* 0x8de2 */
            {8'h00}, /* 0x8de1 */
            {8'h00}, /* 0x8de0 */
            {8'h00}, /* 0x8ddf */
            {8'h00}, /* 0x8dde */
            {8'h00}, /* 0x8ddd */
            {8'h00}, /* 0x8ddc */
            {8'h00}, /* 0x8ddb */
            {8'h00}, /* 0x8dda */
            {8'h00}, /* 0x8dd9 */
            {8'h00}, /* 0x8dd8 */
            {8'h00}, /* 0x8dd7 */
            {8'h00}, /* 0x8dd6 */
            {8'h00}, /* 0x8dd5 */
            {8'h00}, /* 0x8dd4 */
            {8'h00}, /* 0x8dd3 */
            {8'h00}, /* 0x8dd2 */
            {8'h00}, /* 0x8dd1 */
            {8'h00}, /* 0x8dd0 */
            {8'h00}, /* 0x8dcf */
            {8'h00}, /* 0x8dce */
            {8'h00}, /* 0x8dcd */
            {8'h00}, /* 0x8dcc */
            {8'h00}, /* 0x8dcb */
            {8'h00}, /* 0x8dca */
            {8'h00}, /* 0x8dc9 */
            {8'h00}, /* 0x8dc8 */
            {8'h00}, /* 0x8dc7 */
            {8'h00}, /* 0x8dc6 */
            {8'h00}, /* 0x8dc5 */
            {8'h00}, /* 0x8dc4 */
            {8'h00}, /* 0x8dc3 */
            {8'h00}, /* 0x8dc2 */
            {8'h00}, /* 0x8dc1 */
            {8'h00}, /* 0x8dc0 */
            {8'h00}, /* 0x8dbf */
            {8'h00}, /* 0x8dbe */
            {8'h00}, /* 0x8dbd */
            {8'h00}, /* 0x8dbc */
            {8'h00}, /* 0x8dbb */
            {8'h00}, /* 0x8dba */
            {8'h00}, /* 0x8db9 */
            {8'h00}, /* 0x8db8 */
            {8'h00}, /* 0x8db7 */
            {8'h00}, /* 0x8db6 */
            {8'h00}, /* 0x8db5 */
            {8'h00}, /* 0x8db4 */
            {8'h00}, /* 0x8db3 */
            {8'h00}, /* 0x8db2 */
            {8'h00}, /* 0x8db1 */
            {8'h00}, /* 0x8db0 */
            {8'h00}, /* 0x8daf */
            {8'h00}, /* 0x8dae */
            {8'h00}, /* 0x8dad */
            {8'h00}, /* 0x8dac */
            {8'h00}, /* 0x8dab */
            {8'h00}, /* 0x8daa */
            {8'h00}, /* 0x8da9 */
            {8'h00}, /* 0x8da8 */
            {8'h00}, /* 0x8da7 */
            {8'h00}, /* 0x8da6 */
            {8'h00}, /* 0x8da5 */
            {8'h00}, /* 0x8da4 */
            {8'h00}, /* 0x8da3 */
            {8'h00}, /* 0x8da2 */
            {8'h00}, /* 0x8da1 */
            {8'h00}, /* 0x8da0 */
            {8'h00}, /* 0x8d9f */
            {8'h00}, /* 0x8d9e */
            {8'h00}, /* 0x8d9d */
            {8'h00}, /* 0x8d9c */
            {8'h00}, /* 0x8d9b */
            {8'h00}, /* 0x8d9a */
            {8'h00}, /* 0x8d99 */
            {8'h00}, /* 0x8d98 */
            {8'h00}, /* 0x8d97 */
            {8'h00}, /* 0x8d96 */
            {8'h00}, /* 0x8d95 */
            {8'h00}, /* 0x8d94 */
            {8'h00}, /* 0x8d93 */
            {8'h00}, /* 0x8d92 */
            {8'h00}, /* 0x8d91 */
            {8'h00}, /* 0x8d90 */
            {8'h00}, /* 0x8d8f */
            {8'h00}, /* 0x8d8e */
            {8'h00}, /* 0x8d8d */
            {8'h00}, /* 0x8d8c */
            {8'h00}, /* 0x8d8b */
            {8'h00}, /* 0x8d8a */
            {8'h00}, /* 0x8d89 */
            {8'h00}, /* 0x8d88 */
            {8'h00}, /* 0x8d87 */
            {8'h00}, /* 0x8d86 */
            {8'h00}, /* 0x8d85 */
            {8'h00}, /* 0x8d84 */
            {8'h00}, /* 0x8d83 */
            {8'h00}, /* 0x8d82 */
            {8'h00}, /* 0x8d81 */
            {8'h00}, /* 0x8d80 */
            {8'h00}, /* 0x8d7f */
            {8'h00}, /* 0x8d7e */
            {8'h00}, /* 0x8d7d */
            {8'h00}, /* 0x8d7c */
            {8'h00}, /* 0x8d7b */
            {8'h00}, /* 0x8d7a */
            {8'h00}, /* 0x8d79 */
            {8'h00}, /* 0x8d78 */
            {8'h00}, /* 0x8d77 */
            {8'h00}, /* 0x8d76 */
            {8'h00}, /* 0x8d75 */
            {8'h00}, /* 0x8d74 */
            {8'h00}, /* 0x8d73 */
            {8'h00}, /* 0x8d72 */
            {8'h00}, /* 0x8d71 */
            {8'h00}, /* 0x8d70 */
            {8'h00}, /* 0x8d6f */
            {8'h00}, /* 0x8d6e */
            {8'h00}, /* 0x8d6d */
            {8'h00}, /* 0x8d6c */
            {8'h00}, /* 0x8d6b */
            {8'h00}, /* 0x8d6a */
            {8'h00}, /* 0x8d69 */
            {8'h00}, /* 0x8d68 */
            {8'h00}, /* 0x8d67 */
            {8'h00}, /* 0x8d66 */
            {8'h00}, /* 0x8d65 */
            {8'h00}, /* 0x8d64 */
            {8'h00}, /* 0x8d63 */
            {8'h00}, /* 0x8d62 */
            {8'h00}, /* 0x8d61 */
            {8'h00}, /* 0x8d60 */
            {8'h00}, /* 0x8d5f */
            {8'h00}, /* 0x8d5e */
            {8'h00}, /* 0x8d5d */
            {8'h00}, /* 0x8d5c */
            {8'h00}, /* 0x8d5b */
            {8'h00}, /* 0x8d5a */
            {8'h00}, /* 0x8d59 */
            {8'h00}, /* 0x8d58 */
            {8'h00}, /* 0x8d57 */
            {8'h00}, /* 0x8d56 */
            {8'h00}, /* 0x8d55 */
            {8'h00}, /* 0x8d54 */
            {8'h00}, /* 0x8d53 */
            {8'h00}, /* 0x8d52 */
            {8'h00}, /* 0x8d51 */
            {8'h00}, /* 0x8d50 */
            {8'h00}, /* 0x8d4f */
            {8'h00}, /* 0x8d4e */
            {8'h00}, /* 0x8d4d */
            {8'h00}, /* 0x8d4c */
            {8'h00}, /* 0x8d4b */
            {8'h00}, /* 0x8d4a */
            {8'h00}, /* 0x8d49 */
            {8'h00}, /* 0x8d48 */
            {8'h00}, /* 0x8d47 */
            {8'h00}, /* 0x8d46 */
            {8'h00}, /* 0x8d45 */
            {8'h00}, /* 0x8d44 */
            {8'h00}, /* 0x8d43 */
            {8'h00}, /* 0x8d42 */
            {8'h00}, /* 0x8d41 */
            {8'h00}, /* 0x8d40 */
            {8'h00}, /* 0x8d3f */
            {8'h00}, /* 0x8d3e */
            {8'h00}, /* 0x8d3d */
            {8'h00}, /* 0x8d3c */
            {8'h00}, /* 0x8d3b */
            {8'h00}, /* 0x8d3a */
            {8'h00}, /* 0x8d39 */
            {8'h00}, /* 0x8d38 */
            {8'h00}, /* 0x8d37 */
            {8'h00}, /* 0x8d36 */
            {8'h00}, /* 0x8d35 */
            {8'h00}, /* 0x8d34 */
            {8'h00}, /* 0x8d33 */
            {8'h00}, /* 0x8d32 */
            {8'h00}, /* 0x8d31 */
            {8'h00}, /* 0x8d30 */
            {8'h00}, /* 0x8d2f */
            {8'h00}, /* 0x8d2e */
            {8'h00}, /* 0x8d2d */
            {8'h00}, /* 0x8d2c */
            {8'h00}, /* 0x8d2b */
            {8'h00}, /* 0x8d2a */
            {8'h00}, /* 0x8d29 */
            {8'h00}, /* 0x8d28 */
            {8'h00}, /* 0x8d27 */
            {8'h00}, /* 0x8d26 */
            {8'h00}, /* 0x8d25 */
            {8'h00}, /* 0x8d24 */
            {8'h00}, /* 0x8d23 */
            {8'h00}, /* 0x8d22 */
            {8'h00}, /* 0x8d21 */
            {8'h00}, /* 0x8d20 */
            {8'h00}, /* 0x8d1f */
            {8'h00}, /* 0x8d1e */
            {8'h00}, /* 0x8d1d */
            {8'h00}, /* 0x8d1c */
            {8'h00}, /* 0x8d1b */
            {8'h00}, /* 0x8d1a */
            {8'h00}, /* 0x8d19 */
            {8'h00}, /* 0x8d18 */
            {8'h00}, /* 0x8d17 */
            {8'h00}, /* 0x8d16 */
            {8'h00}, /* 0x8d15 */
            {8'h00}, /* 0x8d14 */
            {8'h00}, /* 0x8d13 */
            {8'h00}, /* 0x8d12 */
            {8'h00}, /* 0x8d11 */
            {8'h00}, /* 0x8d10 */
            {8'h00}, /* 0x8d0f */
            {8'h00}, /* 0x8d0e */
            {8'h00}, /* 0x8d0d */
            {8'h00}, /* 0x8d0c */
            {8'h00}, /* 0x8d0b */
            {8'h00}, /* 0x8d0a */
            {8'h00}, /* 0x8d09 */
            {8'h00}, /* 0x8d08 */
            {8'h00}, /* 0x8d07 */
            {8'h00}, /* 0x8d06 */
            {8'h00}, /* 0x8d05 */
            {8'h00}, /* 0x8d04 */
            {8'h00}, /* 0x8d03 */
            {8'h00}, /* 0x8d02 */
            {8'h00}, /* 0x8d01 */
            {8'h00}, /* 0x8d00 */
            {8'h00}, /* 0x8cff */
            {8'h00}, /* 0x8cfe */
            {8'h00}, /* 0x8cfd */
            {8'h00}, /* 0x8cfc */
            {8'h00}, /* 0x8cfb */
            {8'h00}, /* 0x8cfa */
            {8'h00}, /* 0x8cf9 */
            {8'h00}, /* 0x8cf8 */
            {8'h00}, /* 0x8cf7 */
            {8'h00}, /* 0x8cf6 */
            {8'h00}, /* 0x8cf5 */
            {8'h00}, /* 0x8cf4 */
            {8'h00}, /* 0x8cf3 */
            {8'h00}, /* 0x8cf2 */
            {8'h00}, /* 0x8cf1 */
            {8'h00}, /* 0x8cf0 */
            {8'h00}, /* 0x8cef */
            {8'h00}, /* 0x8cee */
            {8'h00}, /* 0x8ced */
            {8'h00}, /* 0x8cec */
            {8'h00}, /* 0x8ceb */
            {8'h00}, /* 0x8cea */
            {8'h00}, /* 0x8ce9 */
            {8'h00}, /* 0x8ce8 */
            {8'h00}, /* 0x8ce7 */
            {8'h00}, /* 0x8ce6 */
            {8'h00}, /* 0x8ce5 */
            {8'h00}, /* 0x8ce4 */
            {8'h00}, /* 0x8ce3 */
            {8'h00}, /* 0x8ce2 */
            {8'h00}, /* 0x8ce1 */
            {8'h00}, /* 0x8ce0 */
            {8'h00}, /* 0x8cdf */
            {8'h00}, /* 0x8cde */
            {8'h00}, /* 0x8cdd */
            {8'h00}, /* 0x8cdc */
            {8'h00}, /* 0x8cdb */
            {8'h00}, /* 0x8cda */
            {8'h00}, /* 0x8cd9 */
            {8'h00}, /* 0x8cd8 */
            {8'h00}, /* 0x8cd7 */
            {8'h00}, /* 0x8cd6 */
            {8'h00}, /* 0x8cd5 */
            {8'h00}, /* 0x8cd4 */
            {8'h00}, /* 0x8cd3 */
            {8'h00}, /* 0x8cd2 */
            {8'h00}, /* 0x8cd1 */
            {8'h00}, /* 0x8cd0 */
            {8'h00}, /* 0x8ccf */
            {8'h00}, /* 0x8cce */
            {8'h00}, /* 0x8ccd */
            {8'h00}, /* 0x8ccc */
            {8'h00}, /* 0x8ccb */
            {8'h00}, /* 0x8cca */
            {8'h00}, /* 0x8cc9 */
            {8'h00}, /* 0x8cc8 */
            {8'h00}, /* 0x8cc7 */
            {8'h00}, /* 0x8cc6 */
            {8'h00}, /* 0x8cc5 */
            {8'h00}, /* 0x8cc4 */
            {8'h00}, /* 0x8cc3 */
            {8'h00}, /* 0x8cc2 */
            {8'h00}, /* 0x8cc1 */
            {8'h00}, /* 0x8cc0 */
            {8'h00}, /* 0x8cbf */
            {8'h00}, /* 0x8cbe */
            {8'h00}, /* 0x8cbd */
            {8'h00}, /* 0x8cbc */
            {8'h00}, /* 0x8cbb */
            {8'h00}, /* 0x8cba */
            {8'h00}, /* 0x8cb9 */
            {8'h00}, /* 0x8cb8 */
            {8'h00}, /* 0x8cb7 */
            {8'h00}, /* 0x8cb6 */
            {8'h00}, /* 0x8cb5 */
            {8'h00}, /* 0x8cb4 */
            {8'h00}, /* 0x8cb3 */
            {8'h00}, /* 0x8cb2 */
            {8'h00}, /* 0x8cb1 */
            {8'h00}, /* 0x8cb0 */
            {8'h00}, /* 0x8caf */
            {8'h00}, /* 0x8cae */
            {8'h00}, /* 0x8cad */
            {8'h00}, /* 0x8cac */
            {8'h00}, /* 0x8cab */
            {8'h00}, /* 0x8caa */
            {8'h00}, /* 0x8ca9 */
            {8'h00}, /* 0x8ca8 */
            {8'h00}, /* 0x8ca7 */
            {8'h00}, /* 0x8ca6 */
            {8'h00}, /* 0x8ca5 */
            {8'h00}, /* 0x8ca4 */
            {8'h00}, /* 0x8ca3 */
            {8'h00}, /* 0x8ca2 */
            {8'h00}, /* 0x8ca1 */
            {8'h00}, /* 0x8ca0 */
            {8'h00}, /* 0x8c9f */
            {8'h00}, /* 0x8c9e */
            {8'h00}, /* 0x8c9d */
            {8'h00}, /* 0x8c9c */
            {8'h00}, /* 0x8c9b */
            {8'h00}, /* 0x8c9a */
            {8'h00}, /* 0x8c99 */
            {8'h00}, /* 0x8c98 */
            {8'h00}, /* 0x8c97 */
            {8'h00}, /* 0x8c96 */
            {8'h00}, /* 0x8c95 */
            {8'h00}, /* 0x8c94 */
            {8'h00}, /* 0x8c93 */
            {8'h00}, /* 0x8c92 */
            {8'h00}, /* 0x8c91 */
            {8'h00}, /* 0x8c90 */
            {8'h00}, /* 0x8c8f */
            {8'h00}, /* 0x8c8e */
            {8'h00}, /* 0x8c8d */
            {8'h00}, /* 0x8c8c */
            {8'h00}, /* 0x8c8b */
            {8'h00}, /* 0x8c8a */
            {8'h00}, /* 0x8c89 */
            {8'h00}, /* 0x8c88 */
            {8'h00}, /* 0x8c87 */
            {8'h00}, /* 0x8c86 */
            {8'h00}, /* 0x8c85 */
            {8'h00}, /* 0x8c84 */
            {8'h00}, /* 0x8c83 */
            {8'h00}, /* 0x8c82 */
            {8'h00}, /* 0x8c81 */
            {8'h00}, /* 0x8c80 */
            {8'h00}, /* 0x8c7f */
            {8'h00}, /* 0x8c7e */
            {8'h00}, /* 0x8c7d */
            {8'h00}, /* 0x8c7c */
            {8'h00}, /* 0x8c7b */
            {8'h00}, /* 0x8c7a */
            {8'h00}, /* 0x8c79 */
            {8'h00}, /* 0x8c78 */
            {8'h00}, /* 0x8c77 */
            {8'h00}, /* 0x8c76 */
            {8'h00}, /* 0x8c75 */
            {8'h00}, /* 0x8c74 */
            {8'h00}, /* 0x8c73 */
            {8'h00}, /* 0x8c72 */
            {8'h00}, /* 0x8c71 */
            {8'h00}, /* 0x8c70 */
            {8'h00}, /* 0x8c6f */
            {8'h00}, /* 0x8c6e */
            {8'h00}, /* 0x8c6d */
            {8'h00}, /* 0x8c6c */
            {8'h00}, /* 0x8c6b */
            {8'h00}, /* 0x8c6a */
            {8'h00}, /* 0x8c69 */
            {8'h00}, /* 0x8c68 */
            {8'h00}, /* 0x8c67 */
            {8'h00}, /* 0x8c66 */
            {8'h00}, /* 0x8c65 */
            {8'h00}, /* 0x8c64 */
            {8'h00}, /* 0x8c63 */
            {8'h00}, /* 0x8c62 */
            {8'h00}, /* 0x8c61 */
            {8'h00}, /* 0x8c60 */
            {8'h00}, /* 0x8c5f */
            {8'h00}, /* 0x8c5e */
            {8'h00}, /* 0x8c5d */
            {8'h00}, /* 0x8c5c */
            {8'h00}, /* 0x8c5b */
            {8'h00}, /* 0x8c5a */
            {8'h00}, /* 0x8c59 */
            {8'h00}, /* 0x8c58 */
            {8'h00}, /* 0x8c57 */
            {8'h00}, /* 0x8c56 */
            {8'h00}, /* 0x8c55 */
            {8'h00}, /* 0x8c54 */
            {8'h00}, /* 0x8c53 */
            {8'h00}, /* 0x8c52 */
            {8'h00}, /* 0x8c51 */
            {8'h00}, /* 0x8c50 */
            {8'h00}, /* 0x8c4f */
            {8'h00}, /* 0x8c4e */
            {8'h00}, /* 0x8c4d */
            {8'h00}, /* 0x8c4c */
            {8'h00}, /* 0x8c4b */
            {8'h00}, /* 0x8c4a */
            {8'h00}, /* 0x8c49 */
            {8'h00}, /* 0x8c48 */
            {8'h00}, /* 0x8c47 */
            {8'h00}, /* 0x8c46 */
            {8'h00}, /* 0x8c45 */
            {8'h00}, /* 0x8c44 */
            {8'h00}, /* 0x8c43 */
            {8'h00}, /* 0x8c42 */
            {8'h00}, /* 0x8c41 */
            {8'h00}, /* 0x8c40 */
            {8'h00}, /* 0x8c3f */
            {8'h00}, /* 0x8c3e */
            {8'h00}, /* 0x8c3d */
            {8'h00}, /* 0x8c3c */
            {8'h00}, /* 0x8c3b */
            {8'h00}, /* 0x8c3a */
            {8'h00}, /* 0x8c39 */
            {8'h00}, /* 0x8c38 */
            {8'h00}, /* 0x8c37 */
            {8'h00}, /* 0x8c36 */
            {8'h00}, /* 0x8c35 */
            {8'h00}, /* 0x8c34 */
            {8'h00}, /* 0x8c33 */
            {8'h00}, /* 0x8c32 */
            {8'h00}, /* 0x8c31 */
            {8'h00}, /* 0x8c30 */
            {8'h00}, /* 0x8c2f */
            {8'h00}, /* 0x8c2e */
            {8'h00}, /* 0x8c2d */
            {8'h00}, /* 0x8c2c */
            {8'h00}, /* 0x8c2b */
            {8'h00}, /* 0x8c2a */
            {8'h00}, /* 0x8c29 */
            {8'h00}, /* 0x8c28 */
            {8'h00}, /* 0x8c27 */
            {8'h00}, /* 0x8c26 */
            {8'h00}, /* 0x8c25 */
            {8'h00}, /* 0x8c24 */
            {8'h00}, /* 0x8c23 */
            {8'h00}, /* 0x8c22 */
            {8'h00}, /* 0x8c21 */
            {8'h00}, /* 0x8c20 */
            {8'h00}, /* 0x8c1f */
            {8'h00}, /* 0x8c1e */
            {8'h00}, /* 0x8c1d */
            {8'h00}, /* 0x8c1c */
            {8'h00}, /* 0x8c1b */
            {8'h00}, /* 0x8c1a */
            {8'h00}, /* 0x8c19 */
            {8'h00}, /* 0x8c18 */
            {8'h00}, /* 0x8c17 */
            {8'h00}, /* 0x8c16 */
            {8'h00}, /* 0x8c15 */
            {8'h00}, /* 0x8c14 */
            {8'h00}, /* 0x8c13 */
            {8'h00}, /* 0x8c12 */
            {8'h00}, /* 0x8c11 */
            {8'h00}, /* 0x8c10 */
            {8'h00}, /* 0x8c0f */
            {8'h00}, /* 0x8c0e */
            {8'h00}, /* 0x8c0d */
            {8'h00}, /* 0x8c0c */
            {8'h00}, /* 0x8c0b */
            {8'h00}, /* 0x8c0a */
            {8'h00}, /* 0x8c09 */
            {8'h00}, /* 0x8c08 */
            {8'h00}, /* 0x8c07 */
            {8'h00}, /* 0x8c06 */
            {8'h00}, /* 0x8c05 */
            {8'h00}, /* 0x8c04 */
            {8'h00}, /* 0x8c03 */
            {8'h00}, /* 0x8c02 */
            {8'h00}, /* 0x8c01 */
            {8'h00}, /* 0x8c00 */
            {8'h00}, /* 0x8bff */
            {8'h00}, /* 0x8bfe */
            {8'h00}, /* 0x8bfd */
            {8'h00}, /* 0x8bfc */
            {8'h00}, /* 0x8bfb */
            {8'h00}, /* 0x8bfa */
            {8'h00}, /* 0x8bf9 */
            {8'h00}, /* 0x8bf8 */
            {8'h00}, /* 0x8bf7 */
            {8'h00}, /* 0x8bf6 */
            {8'h00}, /* 0x8bf5 */
            {8'h00}, /* 0x8bf4 */
            {8'h00}, /* 0x8bf3 */
            {8'h00}, /* 0x8bf2 */
            {8'h00}, /* 0x8bf1 */
            {8'h00}, /* 0x8bf0 */
            {8'h00}, /* 0x8bef */
            {8'h00}, /* 0x8bee */
            {8'h00}, /* 0x8bed */
            {8'h00}, /* 0x8bec */
            {8'h00}, /* 0x8beb */
            {8'h00}, /* 0x8bea */
            {8'h00}, /* 0x8be9 */
            {8'h00}, /* 0x8be8 */
            {8'h00}, /* 0x8be7 */
            {8'h00}, /* 0x8be6 */
            {8'h00}, /* 0x8be5 */
            {8'h00}, /* 0x8be4 */
            {8'h00}, /* 0x8be3 */
            {8'h00}, /* 0x8be2 */
            {8'h00}, /* 0x8be1 */
            {8'h00}, /* 0x8be0 */
            {8'h00}, /* 0x8bdf */
            {8'h00}, /* 0x8bde */
            {8'h00}, /* 0x8bdd */
            {8'h00}, /* 0x8bdc */
            {8'h00}, /* 0x8bdb */
            {8'h00}, /* 0x8bda */
            {8'h00}, /* 0x8bd9 */
            {8'h00}, /* 0x8bd8 */
            {8'h00}, /* 0x8bd7 */
            {8'h00}, /* 0x8bd6 */
            {8'h00}, /* 0x8bd5 */
            {8'h00}, /* 0x8bd4 */
            {8'h00}, /* 0x8bd3 */
            {8'h00}, /* 0x8bd2 */
            {8'h00}, /* 0x8bd1 */
            {8'h00}, /* 0x8bd0 */
            {8'h00}, /* 0x8bcf */
            {8'h00}, /* 0x8bce */
            {8'h00}, /* 0x8bcd */
            {8'h00}, /* 0x8bcc */
            {8'h00}, /* 0x8bcb */
            {8'h00}, /* 0x8bca */
            {8'h00}, /* 0x8bc9 */
            {8'h00}, /* 0x8bc8 */
            {8'h00}, /* 0x8bc7 */
            {8'h00}, /* 0x8bc6 */
            {8'h00}, /* 0x8bc5 */
            {8'h00}, /* 0x8bc4 */
            {8'h00}, /* 0x8bc3 */
            {8'h00}, /* 0x8bc2 */
            {8'h00}, /* 0x8bc1 */
            {8'h00}, /* 0x8bc0 */
            {8'h00}, /* 0x8bbf */
            {8'h00}, /* 0x8bbe */
            {8'h00}, /* 0x8bbd */
            {8'h00}, /* 0x8bbc */
            {8'h00}, /* 0x8bbb */
            {8'h00}, /* 0x8bba */
            {8'h00}, /* 0x8bb9 */
            {8'h00}, /* 0x8bb8 */
            {8'h00}, /* 0x8bb7 */
            {8'h00}, /* 0x8bb6 */
            {8'h00}, /* 0x8bb5 */
            {8'h00}, /* 0x8bb4 */
            {8'h00}, /* 0x8bb3 */
            {8'h00}, /* 0x8bb2 */
            {8'h00}, /* 0x8bb1 */
            {8'h00}, /* 0x8bb0 */
            {8'h00}, /* 0x8baf */
            {8'h00}, /* 0x8bae */
            {8'h00}, /* 0x8bad */
            {8'h00}, /* 0x8bac */
            {8'h00}, /* 0x8bab */
            {8'h00}, /* 0x8baa */
            {8'h00}, /* 0x8ba9 */
            {8'h00}, /* 0x8ba8 */
            {8'h00}, /* 0x8ba7 */
            {8'h00}, /* 0x8ba6 */
            {8'h00}, /* 0x8ba5 */
            {8'h00}, /* 0x8ba4 */
            {8'h00}, /* 0x8ba3 */
            {8'h00}, /* 0x8ba2 */
            {8'h00}, /* 0x8ba1 */
            {8'h00}, /* 0x8ba0 */
            {8'h00}, /* 0x8b9f */
            {8'h00}, /* 0x8b9e */
            {8'h00}, /* 0x8b9d */
            {8'h00}, /* 0x8b9c */
            {8'h00}, /* 0x8b9b */
            {8'h00}, /* 0x8b9a */
            {8'h00}, /* 0x8b99 */
            {8'h00}, /* 0x8b98 */
            {8'h00}, /* 0x8b97 */
            {8'h00}, /* 0x8b96 */
            {8'h00}, /* 0x8b95 */
            {8'h00}, /* 0x8b94 */
            {8'h00}, /* 0x8b93 */
            {8'h00}, /* 0x8b92 */
            {8'h00}, /* 0x8b91 */
            {8'h00}, /* 0x8b90 */
            {8'h00}, /* 0x8b8f */
            {8'h00}, /* 0x8b8e */
            {8'h00}, /* 0x8b8d */
            {8'h00}, /* 0x8b8c */
            {8'h00}, /* 0x8b8b */
            {8'h00}, /* 0x8b8a */
            {8'h00}, /* 0x8b89 */
            {8'h00}, /* 0x8b88 */
            {8'h00}, /* 0x8b87 */
            {8'h00}, /* 0x8b86 */
            {8'h00}, /* 0x8b85 */
            {8'h00}, /* 0x8b84 */
            {8'h00}, /* 0x8b83 */
            {8'h00}, /* 0x8b82 */
            {8'h00}, /* 0x8b81 */
            {8'h00}, /* 0x8b80 */
            {8'h00}, /* 0x8b7f */
            {8'h00}, /* 0x8b7e */
            {8'h00}, /* 0x8b7d */
            {8'h00}, /* 0x8b7c */
            {8'h00}, /* 0x8b7b */
            {8'h00}, /* 0x8b7a */
            {8'h00}, /* 0x8b79 */
            {8'h00}, /* 0x8b78 */
            {8'h00}, /* 0x8b77 */
            {8'h00}, /* 0x8b76 */
            {8'h00}, /* 0x8b75 */
            {8'h00}, /* 0x8b74 */
            {8'h00}, /* 0x8b73 */
            {8'h00}, /* 0x8b72 */
            {8'h00}, /* 0x8b71 */
            {8'h00}, /* 0x8b70 */
            {8'h00}, /* 0x8b6f */
            {8'h00}, /* 0x8b6e */
            {8'h00}, /* 0x8b6d */
            {8'h00}, /* 0x8b6c */
            {8'h00}, /* 0x8b6b */
            {8'h00}, /* 0x8b6a */
            {8'h00}, /* 0x8b69 */
            {8'h00}, /* 0x8b68 */
            {8'h00}, /* 0x8b67 */
            {8'h00}, /* 0x8b66 */
            {8'h00}, /* 0x8b65 */
            {8'h00}, /* 0x8b64 */
            {8'h00}, /* 0x8b63 */
            {8'h00}, /* 0x8b62 */
            {8'h00}, /* 0x8b61 */
            {8'h00}, /* 0x8b60 */
            {8'h00}, /* 0x8b5f */
            {8'h00}, /* 0x8b5e */
            {8'h00}, /* 0x8b5d */
            {8'h00}, /* 0x8b5c */
            {8'h00}, /* 0x8b5b */
            {8'h00}, /* 0x8b5a */
            {8'h00}, /* 0x8b59 */
            {8'h00}, /* 0x8b58 */
            {8'h00}, /* 0x8b57 */
            {8'h00}, /* 0x8b56 */
            {8'h00}, /* 0x8b55 */
            {8'h00}, /* 0x8b54 */
            {8'h00}, /* 0x8b53 */
            {8'h00}, /* 0x8b52 */
            {8'h00}, /* 0x8b51 */
            {8'h00}, /* 0x8b50 */
            {8'h00}, /* 0x8b4f */
            {8'h00}, /* 0x8b4e */
            {8'h00}, /* 0x8b4d */
            {8'h00}, /* 0x8b4c */
            {8'h00}, /* 0x8b4b */
            {8'h00}, /* 0x8b4a */
            {8'h00}, /* 0x8b49 */
            {8'h00}, /* 0x8b48 */
            {8'h00}, /* 0x8b47 */
            {8'h00}, /* 0x8b46 */
            {8'h00}, /* 0x8b45 */
            {8'h00}, /* 0x8b44 */
            {8'h00}, /* 0x8b43 */
            {8'h00}, /* 0x8b42 */
            {8'h00}, /* 0x8b41 */
            {8'h00}, /* 0x8b40 */
            {8'h00}, /* 0x8b3f */
            {8'h00}, /* 0x8b3e */
            {8'h00}, /* 0x8b3d */
            {8'h00}, /* 0x8b3c */
            {8'h00}, /* 0x8b3b */
            {8'h00}, /* 0x8b3a */
            {8'h00}, /* 0x8b39 */
            {8'h00}, /* 0x8b38 */
            {8'h00}, /* 0x8b37 */
            {8'h00}, /* 0x8b36 */
            {8'h00}, /* 0x8b35 */
            {8'h00}, /* 0x8b34 */
            {8'h00}, /* 0x8b33 */
            {8'h00}, /* 0x8b32 */
            {8'h00}, /* 0x8b31 */
            {8'h00}, /* 0x8b30 */
            {8'h00}, /* 0x8b2f */
            {8'h00}, /* 0x8b2e */
            {8'h00}, /* 0x8b2d */
            {8'h00}, /* 0x8b2c */
            {8'h00}, /* 0x8b2b */
            {8'h00}, /* 0x8b2a */
            {8'h00}, /* 0x8b29 */
            {8'h00}, /* 0x8b28 */
            {8'h00}, /* 0x8b27 */
            {8'h00}, /* 0x8b26 */
            {8'h00}, /* 0x8b25 */
            {8'h00}, /* 0x8b24 */
            {8'h00}, /* 0x8b23 */
            {8'h00}, /* 0x8b22 */
            {8'h00}, /* 0x8b21 */
            {8'h00}, /* 0x8b20 */
            {8'h00}, /* 0x8b1f */
            {8'h00}, /* 0x8b1e */
            {8'h00}, /* 0x8b1d */
            {8'h00}, /* 0x8b1c */
            {8'h00}, /* 0x8b1b */
            {8'h00}, /* 0x8b1a */
            {8'h00}, /* 0x8b19 */
            {8'h00}, /* 0x8b18 */
            {8'h00}, /* 0x8b17 */
            {8'h00}, /* 0x8b16 */
            {8'h00}, /* 0x8b15 */
            {8'h00}, /* 0x8b14 */
            {8'h00}, /* 0x8b13 */
            {8'h00}, /* 0x8b12 */
            {8'h00}, /* 0x8b11 */
            {8'h00}, /* 0x8b10 */
            {8'h00}, /* 0x8b0f */
            {8'h00}, /* 0x8b0e */
            {8'h00}, /* 0x8b0d */
            {8'h00}, /* 0x8b0c */
            {8'h00}, /* 0x8b0b */
            {8'h00}, /* 0x8b0a */
            {8'h00}, /* 0x8b09 */
            {8'h00}, /* 0x8b08 */
            {8'h00}, /* 0x8b07 */
            {8'h00}, /* 0x8b06 */
            {8'h00}, /* 0x8b05 */
            {8'h00}, /* 0x8b04 */
            {8'h00}, /* 0x8b03 */
            {8'h00}, /* 0x8b02 */
            {8'h00}, /* 0x8b01 */
            {8'h00}, /* 0x8b00 */
            {8'h00}, /* 0x8aff */
            {8'h00}, /* 0x8afe */
            {8'h00}, /* 0x8afd */
            {8'h00}, /* 0x8afc */
            {8'h00}, /* 0x8afb */
            {8'h00}, /* 0x8afa */
            {8'h00}, /* 0x8af9 */
            {8'h00}, /* 0x8af8 */
            {8'h00}, /* 0x8af7 */
            {8'h00}, /* 0x8af6 */
            {8'h00}, /* 0x8af5 */
            {8'h00}, /* 0x8af4 */
            {8'h00}, /* 0x8af3 */
            {8'h00}, /* 0x8af2 */
            {8'h00}, /* 0x8af1 */
            {8'h00}, /* 0x8af0 */
            {8'h00}, /* 0x8aef */
            {8'h00}, /* 0x8aee */
            {8'h00}, /* 0x8aed */
            {8'h00}, /* 0x8aec */
            {8'h00}, /* 0x8aeb */
            {8'h00}, /* 0x8aea */
            {8'h00}, /* 0x8ae9 */
            {8'h00}, /* 0x8ae8 */
            {8'h00}, /* 0x8ae7 */
            {8'h00}, /* 0x8ae6 */
            {8'h00}, /* 0x8ae5 */
            {8'h00}, /* 0x8ae4 */
            {8'h00}, /* 0x8ae3 */
            {8'h00}, /* 0x8ae2 */
            {8'h00}, /* 0x8ae1 */
            {8'h00}, /* 0x8ae0 */
            {8'h00}, /* 0x8adf */
            {8'h00}, /* 0x8ade */
            {8'h00}, /* 0x8add */
            {8'h00}, /* 0x8adc */
            {8'h00}, /* 0x8adb */
            {8'h00}, /* 0x8ada */
            {8'h00}, /* 0x8ad9 */
            {8'h00}, /* 0x8ad8 */
            {8'h00}, /* 0x8ad7 */
            {8'h00}, /* 0x8ad6 */
            {8'h00}, /* 0x8ad5 */
            {8'h00}, /* 0x8ad4 */
            {8'h00}, /* 0x8ad3 */
            {8'h00}, /* 0x8ad2 */
            {8'h00}, /* 0x8ad1 */
            {8'h00}, /* 0x8ad0 */
            {8'h00}, /* 0x8acf */
            {8'h00}, /* 0x8ace */
            {8'h00}, /* 0x8acd */
            {8'h00}, /* 0x8acc */
            {8'h00}, /* 0x8acb */
            {8'h00}, /* 0x8aca */
            {8'h00}, /* 0x8ac9 */
            {8'h00}, /* 0x8ac8 */
            {8'h00}, /* 0x8ac7 */
            {8'h00}, /* 0x8ac6 */
            {8'h00}, /* 0x8ac5 */
            {8'h00}, /* 0x8ac4 */
            {8'h00}, /* 0x8ac3 */
            {8'h00}, /* 0x8ac2 */
            {8'h00}, /* 0x8ac1 */
            {8'h00}, /* 0x8ac0 */
            {8'h00}, /* 0x8abf */
            {8'h00}, /* 0x8abe */
            {8'h00}, /* 0x8abd */
            {8'h00}, /* 0x8abc */
            {8'h00}, /* 0x8abb */
            {8'h00}, /* 0x8aba */
            {8'h00}, /* 0x8ab9 */
            {8'h00}, /* 0x8ab8 */
            {8'h00}, /* 0x8ab7 */
            {8'h00}, /* 0x8ab6 */
            {8'h00}, /* 0x8ab5 */
            {8'h00}, /* 0x8ab4 */
            {8'h00}, /* 0x8ab3 */
            {8'h00}, /* 0x8ab2 */
            {8'h00}, /* 0x8ab1 */
            {8'h00}, /* 0x8ab0 */
            {8'h00}, /* 0x8aaf */
            {8'h00}, /* 0x8aae */
            {8'h00}, /* 0x8aad */
            {8'h00}, /* 0x8aac */
            {8'h00}, /* 0x8aab */
            {8'h00}, /* 0x8aaa */
            {8'h00}, /* 0x8aa9 */
            {8'h00}, /* 0x8aa8 */
            {8'h00}, /* 0x8aa7 */
            {8'h00}, /* 0x8aa6 */
            {8'h00}, /* 0x8aa5 */
            {8'h00}, /* 0x8aa4 */
            {8'h00}, /* 0x8aa3 */
            {8'h00}, /* 0x8aa2 */
            {8'h00}, /* 0x8aa1 */
            {8'h00}, /* 0x8aa0 */
            {8'h00}, /* 0x8a9f */
            {8'h00}, /* 0x8a9e */
            {8'h00}, /* 0x8a9d */
            {8'h00}, /* 0x8a9c */
            {8'h00}, /* 0x8a9b */
            {8'h00}, /* 0x8a9a */
            {8'h00}, /* 0x8a99 */
            {8'h00}, /* 0x8a98 */
            {8'h00}, /* 0x8a97 */
            {8'h00}, /* 0x8a96 */
            {8'h00}, /* 0x8a95 */
            {8'h00}, /* 0x8a94 */
            {8'h00}, /* 0x8a93 */
            {8'h00}, /* 0x8a92 */
            {8'h00}, /* 0x8a91 */
            {8'h00}, /* 0x8a90 */
            {8'h00}, /* 0x8a8f */
            {8'h00}, /* 0x8a8e */
            {8'h00}, /* 0x8a8d */
            {8'h00}, /* 0x8a8c */
            {8'h00}, /* 0x8a8b */
            {8'h00}, /* 0x8a8a */
            {8'h00}, /* 0x8a89 */
            {8'h00}, /* 0x8a88 */
            {8'h00}, /* 0x8a87 */
            {8'h00}, /* 0x8a86 */
            {8'h00}, /* 0x8a85 */
            {8'h00}, /* 0x8a84 */
            {8'h00}, /* 0x8a83 */
            {8'h00}, /* 0x8a82 */
            {8'h00}, /* 0x8a81 */
            {8'h00}, /* 0x8a80 */
            {8'h00}, /* 0x8a7f */
            {8'h00}, /* 0x8a7e */
            {8'h00}, /* 0x8a7d */
            {8'h00}, /* 0x8a7c */
            {8'h00}, /* 0x8a7b */
            {8'h00}, /* 0x8a7a */
            {8'h00}, /* 0x8a79 */
            {8'h00}, /* 0x8a78 */
            {8'h00}, /* 0x8a77 */
            {8'h00}, /* 0x8a76 */
            {8'h00}, /* 0x8a75 */
            {8'h00}, /* 0x8a74 */
            {8'h00}, /* 0x8a73 */
            {8'h00}, /* 0x8a72 */
            {8'h00}, /* 0x8a71 */
            {8'h00}, /* 0x8a70 */
            {8'h00}, /* 0x8a6f */
            {8'h00}, /* 0x8a6e */
            {8'h00}, /* 0x8a6d */
            {8'h00}, /* 0x8a6c */
            {8'h00}, /* 0x8a6b */
            {8'h00}, /* 0x8a6a */
            {8'h00}, /* 0x8a69 */
            {8'h00}, /* 0x8a68 */
            {8'h00}, /* 0x8a67 */
            {8'h00}, /* 0x8a66 */
            {8'h00}, /* 0x8a65 */
            {8'h00}, /* 0x8a64 */
            {8'h00}, /* 0x8a63 */
            {8'h00}, /* 0x8a62 */
            {8'h00}, /* 0x8a61 */
            {8'h00}, /* 0x8a60 */
            {8'h00}, /* 0x8a5f */
            {8'h00}, /* 0x8a5e */
            {8'h00}, /* 0x8a5d */
            {8'h00}, /* 0x8a5c */
            {8'h00}, /* 0x8a5b */
            {8'h00}, /* 0x8a5a */
            {8'h00}, /* 0x8a59 */
            {8'h00}, /* 0x8a58 */
            {8'h00}, /* 0x8a57 */
            {8'h00}, /* 0x8a56 */
            {8'h00}, /* 0x8a55 */
            {8'h00}, /* 0x8a54 */
            {8'h00}, /* 0x8a53 */
            {8'h00}, /* 0x8a52 */
            {8'h00}, /* 0x8a51 */
            {8'h00}, /* 0x8a50 */
            {8'h00}, /* 0x8a4f */
            {8'h00}, /* 0x8a4e */
            {8'h00}, /* 0x8a4d */
            {8'h00}, /* 0x8a4c */
            {8'h00}, /* 0x8a4b */
            {8'h00}, /* 0x8a4a */
            {8'h00}, /* 0x8a49 */
            {8'h00}, /* 0x8a48 */
            {8'h00}, /* 0x8a47 */
            {8'h00}, /* 0x8a46 */
            {8'h00}, /* 0x8a45 */
            {8'h00}, /* 0x8a44 */
            {8'h00}, /* 0x8a43 */
            {8'h00}, /* 0x8a42 */
            {8'h00}, /* 0x8a41 */
            {8'h00}, /* 0x8a40 */
            {8'h00}, /* 0x8a3f */
            {8'h00}, /* 0x8a3e */
            {8'h00}, /* 0x8a3d */
            {8'h00}, /* 0x8a3c */
            {8'h00}, /* 0x8a3b */
            {8'h00}, /* 0x8a3a */
            {8'h00}, /* 0x8a39 */
            {8'h00}, /* 0x8a38 */
            {8'h00}, /* 0x8a37 */
            {8'h00}, /* 0x8a36 */
            {8'h00}, /* 0x8a35 */
            {8'h00}, /* 0x8a34 */
            {8'h00}, /* 0x8a33 */
            {8'h00}, /* 0x8a32 */
            {8'h00}, /* 0x8a31 */
            {8'h00}, /* 0x8a30 */
            {8'h00}, /* 0x8a2f */
            {8'h00}, /* 0x8a2e */
            {8'h00}, /* 0x8a2d */
            {8'h00}, /* 0x8a2c */
            {8'h00}, /* 0x8a2b */
            {8'h00}, /* 0x8a2a */
            {8'h00}, /* 0x8a29 */
            {8'h00}, /* 0x8a28 */
            {8'h00}, /* 0x8a27 */
            {8'h00}, /* 0x8a26 */
            {8'h00}, /* 0x8a25 */
            {8'h00}, /* 0x8a24 */
            {8'h00}, /* 0x8a23 */
            {8'h00}, /* 0x8a22 */
            {8'h00}, /* 0x8a21 */
            {8'h00}, /* 0x8a20 */
            {8'h00}, /* 0x8a1f */
            {8'h00}, /* 0x8a1e */
            {8'h00}, /* 0x8a1d */
            {8'h00}, /* 0x8a1c */
            {8'h00}, /* 0x8a1b */
            {8'h00}, /* 0x8a1a */
            {8'h00}, /* 0x8a19 */
            {8'h00}, /* 0x8a18 */
            {8'h00}, /* 0x8a17 */
            {8'h00}, /* 0x8a16 */
            {8'h00}, /* 0x8a15 */
            {8'h00}, /* 0x8a14 */
            {8'h00}, /* 0x8a13 */
            {8'h00}, /* 0x8a12 */
            {8'h00}, /* 0x8a11 */
            {8'h00}, /* 0x8a10 */
            {8'h00}, /* 0x8a0f */
            {8'h00}, /* 0x8a0e */
            {8'h00}, /* 0x8a0d */
            {8'h00}, /* 0x8a0c */
            {8'h00}, /* 0x8a0b */
            {8'h00}, /* 0x8a0a */
            {8'h00}, /* 0x8a09 */
            {8'h00}, /* 0x8a08 */
            {8'h00}, /* 0x8a07 */
            {8'h00}, /* 0x8a06 */
            {8'h00}, /* 0x8a05 */
            {8'h00}, /* 0x8a04 */
            {8'h00}, /* 0x8a03 */
            {8'h00}, /* 0x8a02 */
            {8'h00}, /* 0x8a01 */
            {8'h00}, /* 0x8a00 */
            {8'h00}, /* 0x89ff */
            {8'h00}, /* 0x89fe */
            {8'h00}, /* 0x89fd */
            {8'h00}, /* 0x89fc */
            {8'h00}, /* 0x89fb */
            {8'h00}, /* 0x89fa */
            {8'h00}, /* 0x89f9 */
            {8'h00}, /* 0x89f8 */
            {8'h00}, /* 0x89f7 */
            {8'h00}, /* 0x89f6 */
            {8'h00}, /* 0x89f5 */
            {8'h00}, /* 0x89f4 */
            {8'h00}, /* 0x89f3 */
            {8'h00}, /* 0x89f2 */
            {8'h00}, /* 0x89f1 */
            {8'h00}, /* 0x89f0 */
            {8'h00}, /* 0x89ef */
            {8'h00}, /* 0x89ee */
            {8'h00}, /* 0x89ed */
            {8'h00}, /* 0x89ec */
            {8'h00}, /* 0x89eb */
            {8'h00}, /* 0x89ea */
            {8'h00}, /* 0x89e9 */
            {8'h00}, /* 0x89e8 */
            {8'h00}, /* 0x89e7 */
            {8'h00}, /* 0x89e6 */
            {8'h00}, /* 0x89e5 */
            {8'h00}, /* 0x89e4 */
            {8'h00}, /* 0x89e3 */
            {8'h00}, /* 0x89e2 */
            {8'h00}, /* 0x89e1 */
            {8'h00}, /* 0x89e0 */
            {8'h00}, /* 0x89df */
            {8'h00}, /* 0x89de */
            {8'h00}, /* 0x89dd */
            {8'h00}, /* 0x89dc */
            {8'h00}, /* 0x89db */
            {8'h00}, /* 0x89da */
            {8'h00}, /* 0x89d9 */
            {8'h00}, /* 0x89d8 */
            {8'h00}, /* 0x89d7 */
            {8'h00}, /* 0x89d6 */
            {8'h00}, /* 0x89d5 */
            {8'h00}, /* 0x89d4 */
            {8'h00}, /* 0x89d3 */
            {8'h00}, /* 0x89d2 */
            {8'h00}, /* 0x89d1 */
            {8'h00}, /* 0x89d0 */
            {8'h00}, /* 0x89cf */
            {8'h00}, /* 0x89ce */
            {8'h00}, /* 0x89cd */
            {8'h00}, /* 0x89cc */
            {8'h00}, /* 0x89cb */
            {8'h00}, /* 0x89ca */
            {8'h00}, /* 0x89c9 */
            {8'h00}, /* 0x89c8 */
            {8'h00}, /* 0x89c7 */
            {8'h00}, /* 0x89c6 */
            {8'h00}, /* 0x89c5 */
            {8'h00}, /* 0x89c4 */
            {8'h00}, /* 0x89c3 */
            {8'h00}, /* 0x89c2 */
            {8'h00}, /* 0x89c1 */
            {8'h00}, /* 0x89c0 */
            {8'h00}, /* 0x89bf */
            {8'h00}, /* 0x89be */
            {8'h00}, /* 0x89bd */
            {8'h00}, /* 0x89bc */
            {8'h00}, /* 0x89bb */
            {8'h00}, /* 0x89ba */
            {8'h00}, /* 0x89b9 */
            {8'h00}, /* 0x89b8 */
            {8'h00}, /* 0x89b7 */
            {8'h00}, /* 0x89b6 */
            {8'h00}, /* 0x89b5 */
            {8'h00}, /* 0x89b4 */
            {8'h00}, /* 0x89b3 */
            {8'h00}, /* 0x89b2 */
            {8'h00}, /* 0x89b1 */
            {8'h00}, /* 0x89b0 */
            {8'h00}, /* 0x89af */
            {8'h00}, /* 0x89ae */
            {8'h00}, /* 0x89ad */
            {8'h00}, /* 0x89ac */
            {8'h00}, /* 0x89ab */
            {8'h00}, /* 0x89aa */
            {8'h00}, /* 0x89a9 */
            {8'h00}, /* 0x89a8 */
            {8'h00}, /* 0x89a7 */
            {8'h00}, /* 0x89a6 */
            {8'h00}, /* 0x89a5 */
            {8'h00}, /* 0x89a4 */
            {8'h00}, /* 0x89a3 */
            {8'h00}, /* 0x89a2 */
            {8'h00}, /* 0x89a1 */
            {8'h00}, /* 0x89a0 */
            {8'h00}, /* 0x899f */
            {8'h00}, /* 0x899e */
            {8'h00}, /* 0x899d */
            {8'h00}, /* 0x899c */
            {8'h00}, /* 0x899b */
            {8'h00}, /* 0x899a */
            {8'h00}, /* 0x8999 */
            {8'h00}, /* 0x8998 */
            {8'h00}, /* 0x8997 */
            {8'h00}, /* 0x8996 */
            {8'h00}, /* 0x8995 */
            {8'h00}, /* 0x8994 */
            {8'h00}, /* 0x8993 */
            {8'h00}, /* 0x8992 */
            {8'h00}, /* 0x8991 */
            {8'h00}, /* 0x8990 */
            {8'h00}, /* 0x898f */
            {8'h00}, /* 0x898e */
            {8'h00}, /* 0x898d */
            {8'h00}, /* 0x898c */
            {8'h00}, /* 0x898b */
            {8'h00}, /* 0x898a */
            {8'h00}, /* 0x8989 */
            {8'h00}, /* 0x8988 */
            {8'h00}, /* 0x8987 */
            {8'h00}, /* 0x8986 */
            {8'h00}, /* 0x8985 */
            {8'h00}, /* 0x8984 */
            {8'h00}, /* 0x8983 */
            {8'h00}, /* 0x8982 */
            {8'h00}, /* 0x8981 */
            {8'h00}, /* 0x8980 */
            {8'h00}, /* 0x897f */
            {8'h00}, /* 0x897e */
            {8'h00}, /* 0x897d */
            {8'h00}, /* 0x897c */
            {8'h00}, /* 0x897b */
            {8'h00}, /* 0x897a */
            {8'h00}, /* 0x8979 */
            {8'h00}, /* 0x8978 */
            {8'h00}, /* 0x8977 */
            {8'h00}, /* 0x8976 */
            {8'h00}, /* 0x8975 */
            {8'h00}, /* 0x8974 */
            {8'h00}, /* 0x8973 */
            {8'h00}, /* 0x8972 */
            {8'h00}, /* 0x8971 */
            {8'h00}, /* 0x8970 */
            {8'h00}, /* 0x896f */
            {8'h00}, /* 0x896e */
            {8'h00}, /* 0x896d */
            {8'h00}, /* 0x896c */
            {8'h00}, /* 0x896b */
            {8'h00}, /* 0x896a */
            {8'h00}, /* 0x8969 */
            {8'h00}, /* 0x8968 */
            {8'h00}, /* 0x8967 */
            {8'h00}, /* 0x8966 */
            {8'h00}, /* 0x8965 */
            {8'h00}, /* 0x8964 */
            {8'h00}, /* 0x8963 */
            {8'h00}, /* 0x8962 */
            {8'h00}, /* 0x8961 */
            {8'h00}, /* 0x8960 */
            {8'h00}, /* 0x895f */
            {8'h00}, /* 0x895e */
            {8'h00}, /* 0x895d */
            {8'h00}, /* 0x895c */
            {8'h00}, /* 0x895b */
            {8'h00}, /* 0x895a */
            {8'h00}, /* 0x8959 */
            {8'h00}, /* 0x8958 */
            {8'h00}, /* 0x8957 */
            {8'h00}, /* 0x8956 */
            {8'h00}, /* 0x8955 */
            {8'h00}, /* 0x8954 */
            {8'h00}, /* 0x8953 */
            {8'h00}, /* 0x8952 */
            {8'h00}, /* 0x8951 */
            {8'h00}, /* 0x8950 */
            {8'h00}, /* 0x894f */
            {8'h00}, /* 0x894e */
            {8'h00}, /* 0x894d */
            {8'h00}, /* 0x894c */
            {8'h00}, /* 0x894b */
            {8'h00}, /* 0x894a */
            {8'h00}, /* 0x8949 */
            {8'h00}, /* 0x8948 */
            {8'h00}, /* 0x8947 */
            {8'h00}, /* 0x8946 */
            {8'h00}, /* 0x8945 */
            {8'h00}, /* 0x8944 */
            {8'h00}, /* 0x8943 */
            {8'h00}, /* 0x8942 */
            {8'h00}, /* 0x8941 */
            {8'h00}, /* 0x8940 */
            {8'h00}, /* 0x893f */
            {8'h00}, /* 0x893e */
            {8'h00}, /* 0x893d */
            {8'h00}, /* 0x893c */
            {8'h00}, /* 0x893b */
            {8'h00}, /* 0x893a */
            {8'h00}, /* 0x8939 */
            {8'h00}, /* 0x8938 */
            {8'h00}, /* 0x8937 */
            {8'h00}, /* 0x8936 */
            {8'h00}, /* 0x8935 */
            {8'h00}, /* 0x8934 */
            {8'h00}, /* 0x8933 */
            {8'h00}, /* 0x8932 */
            {8'h00}, /* 0x8931 */
            {8'h00}, /* 0x8930 */
            {8'h00}, /* 0x892f */
            {8'h00}, /* 0x892e */
            {8'h00}, /* 0x892d */
            {8'h00}, /* 0x892c */
            {8'h00}, /* 0x892b */
            {8'h00}, /* 0x892a */
            {8'h00}, /* 0x8929 */
            {8'h00}, /* 0x8928 */
            {8'h00}, /* 0x8927 */
            {8'h00}, /* 0x8926 */
            {8'h00}, /* 0x8925 */
            {8'h00}, /* 0x8924 */
            {8'h00}, /* 0x8923 */
            {8'h00}, /* 0x8922 */
            {8'h00}, /* 0x8921 */
            {8'h00}, /* 0x8920 */
            {8'h00}, /* 0x891f */
            {8'h00}, /* 0x891e */
            {8'h00}, /* 0x891d */
            {8'h00}, /* 0x891c */
            {8'h00}, /* 0x891b */
            {8'h00}, /* 0x891a */
            {8'h00}, /* 0x8919 */
            {8'h00}, /* 0x8918 */
            {8'h00}, /* 0x8917 */
            {8'h00}, /* 0x8916 */
            {8'h00}, /* 0x8915 */
            {8'h00}, /* 0x8914 */
            {8'h00}, /* 0x8913 */
            {8'h00}, /* 0x8912 */
            {8'h00}, /* 0x8911 */
            {8'h00}, /* 0x8910 */
            {8'h00}, /* 0x890f */
            {8'h00}, /* 0x890e */
            {8'h00}, /* 0x890d */
            {8'h00}, /* 0x890c */
            {8'h00}, /* 0x890b */
            {8'h00}, /* 0x890a */
            {8'h00}, /* 0x8909 */
            {8'h00}, /* 0x8908 */
            {8'h00}, /* 0x8907 */
            {8'h00}, /* 0x8906 */
            {8'h00}, /* 0x8905 */
            {8'h00}, /* 0x8904 */
            {8'h00}, /* 0x8903 */
            {8'h00}, /* 0x8902 */
            {8'h00}, /* 0x8901 */
            {8'h00}, /* 0x8900 */
            {8'h00}, /* 0x88ff */
            {8'h00}, /* 0x88fe */
            {8'h00}, /* 0x88fd */
            {8'h00}, /* 0x88fc */
            {8'h00}, /* 0x88fb */
            {8'h00}, /* 0x88fa */
            {8'h00}, /* 0x88f9 */
            {8'h00}, /* 0x88f8 */
            {8'h00}, /* 0x88f7 */
            {8'h00}, /* 0x88f6 */
            {8'h00}, /* 0x88f5 */
            {8'h00}, /* 0x88f4 */
            {8'h00}, /* 0x88f3 */
            {8'h00}, /* 0x88f2 */
            {8'h00}, /* 0x88f1 */
            {8'h00}, /* 0x88f0 */
            {8'h00}, /* 0x88ef */
            {8'h00}, /* 0x88ee */
            {8'h00}, /* 0x88ed */
            {8'h00}, /* 0x88ec */
            {8'h00}, /* 0x88eb */
            {8'h00}, /* 0x88ea */
            {8'h00}, /* 0x88e9 */
            {8'h00}, /* 0x88e8 */
            {8'h00}, /* 0x88e7 */
            {8'h00}, /* 0x88e6 */
            {8'h00}, /* 0x88e5 */
            {8'h00}, /* 0x88e4 */
            {8'h00}, /* 0x88e3 */
            {8'h00}, /* 0x88e2 */
            {8'h00}, /* 0x88e1 */
            {8'h00}, /* 0x88e0 */
            {8'h00}, /* 0x88df */
            {8'h00}, /* 0x88de */
            {8'h00}, /* 0x88dd */
            {8'h00}, /* 0x88dc */
            {8'h00}, /* 0x88db */
            {8'h00}, /* 0x88da */
            {8'h00}, /* 0x88d9 */
            {8'h00}, /* 0x88d8 */
            {8'h00}, /* 0x88d7 */
            {8'h00}, /* 0x88d6 */
            {8'h00}, /* 0x88d5 */
            {8'h00}, /* 0x88d4 */
            {8'h00}, /* 0x88d3 */
            {8'h00}, /* 0x88d2 */
            {8'h00}, /* 0x88d1 */
            {8'h00}, /* 0x88d0 */
            {8'h00}, /* 0x88cf */
            {8'h00}, /* 0x88ce */
            {8'h00}, /* 0x88cd */
            {8'h00}, /* 0x88cc */
            {8'h00}, /* 0x88cb */
            {8'h00}, /* 0x88ca */
            {8'h00}, /* 0x88c9 */
            {8'h00}, /* 0x88c8 */
            {8'h00}, /* 0x88c7 */
            {8'h00}, /* 0x88c6 */
            {8'h00}, /* 0x88c5 */
            {8'h00}, /* 0x88c4 */
            {8'h00}, /* 0x88c3 */
            {8'h00}, /* 0x88c2 */
            {8'h00}, /* 0x88c1 */
            {8'h00}, /* 0x88c0 */
            {8'h00}, /* 0x88bf */
            {8'h00}, /* 0x88be */
            {8'h00}, /* 0x88bd */
            {8'h00}, /* 0x88bc */
            {8'h00}, /* 0x88bb */
            {8'h00}, /* 0x88ba */
            {8'h00}, /* 0x88b9 */
            {8'h00}, /* 0x88b8 */
            {8'h00}, /* 0x88b7 */
            {8'h00}, /* 0x88b6 */
            {8'h00}, /* 0x88b5 */
            {8'h00}, /* 0x88b4 */
            {8'h00}, /* 0x88b3 */
            {8'h00}, /* 0x88b2 */
            {8'h00}, /* 0x88b1 */
            {8'h00}, /* 0x88b0 */
            {8'h00}, /* 0x88af */
            {8'h00}, /* 0x88ae */
            {8'h00}, /* 0x88ad */
            {8'h00}, /* 0x88ac */
            {8'h00}, /* 0x88ab */
            {8'h00}, /* 0x88aa */
            {8'h00}, /* 0x88a9 */
            {8'h00}, /* 0x88a8 */
            {8'h00}, /* 0x88a7 */
            {8'h00}, /* 0x88a6 */
            {8'h00}, /* 0x88a5 */
            {8'h00}, /* 0x88a4 */
            {8'h00}, /* 0x88a3 */
            {8'h00}, /* 0x88a2 */
            {8'h00}, /* 0x88a1 */
            {8'h00}, /* 0x88a0 */
            {8'h00}, /* 0x889f */
            {8'h00}, /* 0x889e */
            {8'h00}, /* 0x889d */
            {8'h00}, /* 0x889c */
            {8'h00}, /* 0x889b */
            {8'h00}, /* 0x889a */
            {8'h00}, /* 0x8899 */
            {8'h00}, /* 0x8898 */
            {8'h00}, /* 0x8897 */
            {8'h00}, /* 0x8896 */
            {8'h00}, /* 0x8895 */
            {8'h00}, /* 0x8894 */
            {8'h00}, /* 0x8893 */
            {8'h00}, /* 0x8892 */
            {8'h00}, /* 0x8891 */
            {8'h00}, /* 0x8890 */
            {8'h00}, /* 0x888f */
            {8'h00}, /* 0x888e */
            {8'h00}, /* 0x888d */
            {8'h00}, /* 0x888c */
            {8'h00}, /* 0x888b */
            {8'h00}, /* 0x888a */
            {8'h00}, /* 0x8889 */
            {8'h00}, /* 0x8888 */
            {8'h00}, /* 0x8887 */
            {8'h00}, /* 0x8886 */
            {8'h00}, /* 0x8885 */
            {8'h00}, /* 0x8884 */
            {8'h00}, /* 0x8883 */
            {8'h00}, /* 0x8882 */
            {8'h00}, /* 0x8881 */
            {8'h00}, /* 0x8880 */
            {8'h00}, /* 0x887f */
            {8'h00}, /* 0x887e */
            {8'h00}, /* 0x887d */
            {8'h00}, /* 0x887c */
            {8'h00}, /* 0x887b */
            {8'h00}, /* 0x887a */
            {8'h00}, /* 0x8879 */
            {8'h00}, /* 0x8878 */
            {8'h00}, /* 0x8877 */
            {8'h00}, /* 0x8876 */
            {8'h00}, /* 0x8875 */
            {8'h00}, /* 0x8874 */
            {8'h00}, /* 0x8873 */
            {8'h00}, /* 0x8872 */
            {8'h00}, /* 0x8871 */
            {8'h00}, /* 0x8870 */
            {8'h00}, /* 0x886f */
            {8'h00}, /* 0x886e */
            {8'h00}, /* 0x886d */
            {8'h00}, /* 0x886c */
            {8'h00}, /* 0x886b */
            {8'h00}, /* 0x886a */
            {8'h00}, /* 0x8869 */
            {8'h00}, /* 0x8868 */
            {8'h00}, /* 0x8867 */
            {8'h00}, /* 0x8866 */
            {8'h00}, /* 0x8865 */
            {8'h00}, /* 0x8864 */
            {8'h00}, /* 0x8863 */
            {8'h00}, /* 0x8862 */
            {8'h00}, /* 0x8861 */
            {8'h00}, /* 0x8860 */
            {8'h00}, /* 0x885f */
            {8'h00}, /* 0x885e */
            {8'h00}, /* 0x885d */
            {8'h00}, /* 0x885c */
            {8'h00}, /* 0x885b */
            {8'h00}, /* 0x885a */
            {8'h00}, /* 0x8859 */
            {8'h00}, /* 0x8858 */
            {8'h00}, /* 0x8857 */
            {8'h00}, /* 0x8856 */
            {8'h00}, /* 0x8855 */
            {8'h00}, /* 0x8854 */
            {8'h00}, /* 0x8853 */
            {8'h00}, /* 0x8852 */
            {8'h00}, /* 0x8851 */
            {8'h00}, /* 0x8850 */
            {8'h00}, /* 0x884f */
            {8'h00}, /* 0x884e */
            {8'h00}, /* 0x884d */
            {8'h00}, /* 0x884c */
            {8'h00}, /* 0x884b */
            {8'h00}, /* 0x884a */
            {8'h00}, /* 0x8849 */
            {8'h00}, /* 0x8848 */
            {8'h00}, /* 0x8847 */
            {8'h00}, /* 0x8846 */
            {8'h00}, /* 0x8845 */
            {8'h00}, /* 0x8844 */
            {8'h00}, /* 0x8843 */
            {8'h00}, /* 0x8842 */
            {8'h00}, /* 0x8841 */
            {8'h00}, /* 0x8840 */
            {8'h00}, /* 0x883f */
            {8'h00}, /* 0x883e */
            {8'h00}, /* 0x883d */
            {8'h00}, /* 0x883c */
            {8'h00}, /* 0x883b */
            {8'h00}, /* 0x883a */
            {8'h00}, /* 0x8839 */
            {8'h00}, /* 0x8838 */
            {8'h00}, /* 0x8837 */
            {8'h00}, /* 0x8836 */
            {8'h00}, /* 0x8835 */
            {8'h00}, /* 0x8834 */
            {8'h00}, /* 0x8833 */
            {8'h00}, /* 0x8832 */
            {8'h00}, /* 0x8831 */
            {8'h00}, /* 0x8830 */
            {8'h00}, /* 0x882f */
            {8'h00}, /* 0x882e */
            {8'h00}, /* 0x882d */
            {8'h00}, /* 0x882c */
            {8'h00}, /* 0x882b */
            {8'h00}, /* 0x882a */
            {8'h00}, /* 0x8829 */
            {8'h00}, /* 0x8828 */
            {8'h00}, /* 0x8827 */
            {8'h00}, /* 0x8826 */
            {8'h00}, /* 0x8825 */
            {8'h00}, /* 0x8824 */
            {8'h00}, /* 0x8823 */
            {8'h00}, /* 0x8822 */
            {8'h00}, /* 0x8821 */
            {8'h00}, /* 0x8820 */
            {8'h00}, /* 0x881f */
            {8'h00}, /* 0x881e */
            {8'h00}, /* 0x881d */
            {8'h00}, /* 0x881c */
            {8'h00}, /* 0x881b */
            {8'h00}, /* 0x881a */
            {8'h00}, /* 0x8819 */
            {8'h00}, /* 0x8818 */
            {8'h00}, /* 0x8817 */
            {8'h00}, /* 0x8816 */
            {8'h00}, /* 0x8815 */
            {8'h00}, /* 0x8814 */
            {8'h00}, /* 0x8813 */
            {8'h00}, /* 0x8812 */
            {8'h00}, /* 0x8811 */
            {8'h00}, /* 0x8810 */
            {8'h00}, /* 0x880f */
            {8'h00}, /* 0x880e */
            {8'h00}, /* 0x880d */
            {8'h00}, /* 0x880c */
            {8'h00}, /* 0x880b */
            {8'h00}, /* 0x880a */
            {8'h00}, /* 0x8809 */
            {8'h00}, /* 0x8808 */
            {8'h00}, /* 0x8807 */
            {8'h00}, /* 0x8806 */
            {8'h00}, /* 0x8805 */
            {8'h00}, /* 0x8804 */
            {8'h00}, /* 0x8803 */
            {8'h00}, /* 0x8802 */
            {8'h00}, /* 0x8801 */
            {8'h00}, /* 0x8800 */
            {8'h00}, /* 0x87ff */
            {8'h00}, /* 0x87fe */
            {8'h00}, /* 0x87fd */
            {8'h00}, /* 0x87fc */
            {8'h00}, /* 0x87fb */
            {8'h00}, /* 0x87fa */
            {8'h00}, /* 0x87f9 */
            {8'h00}, /* 0x87f8 */
            {8'h00}, /* 0x87f7 */
            {8'h00}, /* 0x87f6 */
            {8'h00}, /* 0x87f5 */
            {8'h00}, /* 0x87f4 */
            {8'h00}, /* 0x87f3 */
            {8'h00}, /* 0x87f2 */
            {8'h00}, /* 0x87f1 */
            {8'h00}, /* 0x87f0 */
            {8'h00}, /* 0x87ef */
            {8'h00}, /* 0x87ee */
            {8'h00}, /* 0x87ed */
            {8'h00}, /* 0x87ec */
            {8'h00}, /* 0x87eb */
            {8'h00}, /* 0x87ea */
            {8'h00}, /* 0x87e9 */
            {8'h00}, /* 0x87e8 */
            {8'h00}, /* 0x87e7 */
            {8'h00}, /* 0x87e6 */
            {8'h00}, /* 0x87e5 */
            {8'h00}, /* 0x87e4 */
            {8'h00}, /* 0x87e3 */
            {8'h00}, /* 0x87e2 */
            {8'h00}, /* 0x87e1 */
            {8'h00}, /* 0x87e0 */
            {8'h00}, /* 0x87df */
            {8'h00}, /* 0x87de */
            {8'h00}, /* 0x87dd */
            {8'h00}, /* 0x87dc */
            {8'h00}, /* 0x87db */
            {8'h00}, /* 0x87da */
            {8'h00}, /* 0x87d9 */
            {8'h00}, /* 0x87d8 */
            {8'h00}, /* 0x87d7 */
            {8'h00}, /* 0x87d6 */
            {8'h00}, /* 0x87d5 */
            {8'h00}, /* 0x87d4 */
            {8'h00}, /* 0x87d3 */
            {8'h00}, /* 0x87d2 */
            {8'h00}, /* 0x87d1 */
            {8'h00}, /* 0x87d0 */
            {8'h00}, /* 0x87cf */
            {8'h00}, /* 0x87ce */
            {8'h00}, /* 0x87cd */
            {8'h00}, /* 0x87cc */
            {8'h00}, /* 0x87cb */
            {8'h00}, /* 0x87ca */
            {8'h00}, /* 0x87c9 */
            {8'h00}, /* 0x87c8 */
            {8'h00}, /* 0x87c7 */
            {8'h00}, /* 0x87c6 */
            {8'h00}, /* 0x87c5 */
            {8'h00}, /* 0x87c4 */
            {8'h00}, /* 0x87c3 */
            {8'h00}, /* 0x87c2 */
            {8'h00}, /* 0x87c1 */
            {8'h00}, /* 0x87c0 */
            {8'h00}, /* 0x87bf */
            {8'h00}, /* 0x87be */
            {8'h00}, /* 0x87bd */
            {8'h00}, /* 0x87bc */
            {8'h00}, /* 0x87bb */
            {8'h00}, /* 0x87ba */
            {8'h00}, /* 0x87b9 */
            {8'h00}, /* 0x87b8 */
            {8'h00}, /* 0x87b7 */
            {8'h00}, /* 0x87b6 */
            {8'h00}, /* 0x87b5 */
            {8'h00}, /* 0x87b4 */
            {8'h00}, /* 0x87b3 */
            {8'h00}, /* 0x87b2 */
            {8'h00}, /* 0x87b1 */
            {8'h00}, /* 0x87b0 */
            {8'h00}, /* 0x87af */
            {8'h00}, /* 0x87ae */
            {8'h00}, /* 0x87ad */
            {8'h00}, /* 0x87ac */
            {8'h00}, /* 0x87ab */
            {8'h00}, /* 0x87aa */
            {8'h00}, /* 0x87a9 */
            {8'h00}, /* 0x87a8 */
            {8'h00}, /* 0x87a7 */
            {8'h00}, /* 0x87a6 */
            {8'h00}, /* 0x87a5 */
            {8'h00}, /* 0x87a4 */
            {8'h00}, /* 0x87a3 */
            {8'h00}, /* 0x87a2 */
            {8'h00}, /* 0x87a1 */
            {8'h00}, /* 0x87a0 */
            {8'h00}, /* 0x879f */
            {8'h00}, /* 0x879e */
            {8'h00}, /* 0x879d */
            {8'h00}, /* 0x879c */
            {8'h00}, /* 0x879b */
            {8'h00}, /* 0x879a */
            {8'h00}, /* 0x8799 */
            {8'h00}, /* 0x8798 */
            {8'h00}, /* 0x8797 */
            {8'h00}, /* 0x8796 */
            {8'h00}, /* 0x8795 */
            {8'h00}, /* 0x8794 */
            {8'h00}, /* 0x8793 */
            {8'h00}, /* 0x8792 */
            {8'h00}, /* 0x8791 */
            {8'h00}, /* 0x8790 */
            {8'h00}, /* 0x878f */
            {8'h00}, /* 0x878e */
            {8'h00}, /* 0x878d */
            {8'h00}, /* 0x878c */
            {8'h00}, /* 0x878b */
            {8'h00}, /* 0x878a */
            {8'h00}, /* 0x8789 */
            {8'h00}, /* 0x8788 */
            {8'h00}, /* 0x8787 */
            {8'h00}, /* 0x8786 */
            {8'h00}, /* 0x8785 */
            {8'h00}, /* 0x8784 */
            {8'h00}, /* 0x8783 */
            {8'h00}, /* 0x8782 */
            {8'h00}, /* 0x8781 */
            {8'h00}, /* 0x8780 */
            {8'h00}, /* 0x877f */
            {8'h00}, /* 0x877e */
            {8'h00}, /* 0x877d */
            {8'h00}, /* 0x877c */
            {8'h00}, /* 0x877b */
            {8'h00}, /* 0x877a */
            {8'h00}, /* 0x8779 */
            {8'h00}, /* 0x8778 */
            {8'h00}, /* 0x8777 */
            {8'h00}, /* 0x8776 */
            {8'h00}, /* 0x8775 */
            {8'h00}, /* 0x8774 */
            {8'h00}, /* 0x8773 */
            {8'h00}, /* 0x8772 */
            {8'h00}, /* 0x8771 */
            {8'h00}, /* 0x8770 */
            {8'h00}, /* 0x876f */
            {8'h00}, /* 0x876e */
            {8'h00}, /* 0x876d */
            {8'h00}, /* 0x876c */
            {8'h00}, /* 0x876b */
            {8'h00}, /* 0x876a */
            {8'h00}, /* 0x8769 */
            {8'h00}, /* 0x8768 */
            {8'h00}, /* 0x8767 */
            {8'h00}, /* 0x8766 */
            {8'h00}, /* 0x8765 */
            {8'h00}, /* 0x8764 */
            {8'h00}, /* 0x8763 */
            {8'h00}, /* 0x8762 */
            {8'h00}, /* 0x8761 */
            {8'h00}, /* 0x8760 */
            {8'h00}, /* 0x875f */
            {8'h00}, /* 0x875e */
            {8'h00}, /* 0x875d */
            {8'h00}, /* 0x875c */
            {8'h00}, /* 0x875b */
            {8'h00}, /* 0x875a */
            {8'h00}, /* 0x8759 */
            {8'h00}, /* 0x8758 */
            {8'h00}, /* 0x8757 */
            {8'h00}, /* 0x8756 */
            {8'h00}, /* 0x8755 */
            {8'h00}, /* 0x8754 */
            {8'h00}, /* 0x8753 */
            {8'h00}, /* 0x8752 */
            {8'h00}, /* 0x8751 */
            {8'h00}, /* 0x8750 */
            {8'h00}, /* 0x874f */
            {8'h00}, /* 0x874e */
            {8'h00}, /* 0x874d */
            {8'h00}, /* 0x874c */
            {8'h00}, /* 0x874b */
            {8'h00}, /* 0x874a */
            {8'h00}, /* 0x8749 */
            {8'h00}, /* 0x8748 */
            {8'h00}, /* 0x8747 */
            {8'h00}, /* 0x8746 */
            {8'h00}, /* 0x8745 */
            {8'h00}, /* 0x8744 */
            {8'h00}, /* 0x8743 */
            {8'h00}, /* 0x8742 */
            {8'h00}, /* 0x8741 */
            {8'h00}, /* 0x8740 */
            {8'h00}, /* 0x873f */
            {8'h00}, /* 0x873e */
            {8'h00}, /* 0x873d */
            {8'h00}, /* 0x873c */
            {8'h00}, /* 0x873b */
            {8'h00}, /* 0x873a */
            {8'h00}, /* 0x8739 */
            {8'h00}, /* 0x8738 */
            {8'h00}, /* 0x8737 */
            {8'h00}, /* 0x8736 */
            {8'h00}, /* 0x8735 */
            {8'h00}, /* 0x8734 */
            {8'h00}, /* 0x8733 */
            {8'h00}, /* 0x8732 */
            {8'h00}, /* 0x8731 */
            {8'h00}, /* 0x8730 */
            {8'h00}, /* 0x872f */
            {8'h00}, /* 0x872e */
            {8'h00}, /* 0x872d */
            {8'h00}, /* 0x872c */
            {8'h00}, /* 0x872b */
            {8'h00}, /* 0x872a */
            {8'h00}, /* 0x8729 */
            {8'h00}, /* 0x8728 */
            {8'h00}, /* 0x8727 */
            {8'h00}, /* 0x8726 */
            {8'h00}, /* 0x8725 */
            {8'h00}, /* 0x8724 */
            {8'h00}, /* 0x8723 */
            {8'h00}, /* 0x8722 */
            {8'h00}, /* 0x8721 */
            {8'h00}, /* 0x8720 */
            {8'h00}, /* 0x871f */
            {8'h00}, /* 0x871e */
            {8'h00}, /* 0x871d */
            {8'h00}, /* 0x871c */
            {8'h00}, /* 0x871b */
            {8'h00}, /* 0x871a */
            {8'h00}, /* 0x8719 */
            {8'h00}, /* 0x8718 */
            {8'h00}, /* 0x8717 */
            {8'h00}, /* 0x8716 */
            {8'h00}, /* 0x8715 */
            {8'h00}, /* 0x8714 */
            {8'h00}, /* 0x8713 */
            {8'h00}, /* 0x8712 */
            {8'h00}, /* 0x8711 */
            {8'h00}, /* 0x8710 */
            {8'h00}, /* 0x870f */
            {8'h00}, /* 0x870e */
            {8'h00}, /* 0x870d */
            {8'h00}, /* 0x870c */
            {8'h00}, /* 0x870b */
            {8'h00}, /* 0x870a */
            {8'h00}, /* 0x8709 */
            {8'h00}, /* 0x8708 */
            {8'h00}, /* 0x8707 */
            {8'h00}, /* 0x8706 */
            {8'h00}, /* 0x8705 */
            {8'h00}, /* 0x8704 */
            {8'h00}, /* 0x8703 */
            {8'h00}, /* 0x8702 */
            {8'h00}, /* 0x8701 */
            {8'h00}, /* 0x8700 */
            {8'h00}, /* 0x86ff */
            {8'h00}, /* 0x86fe */
            {8'h00}, /* 0x86fd */
            {8'h00}, /* 0x86fc */
            {8'h00}, /* 0x86fb */
            {8'h00}, /* 0x86fa */
            {8'h00}, /* 0x86f9 */
            {8'h00}, /* 0x86f8 */
            {8'h00}, /* 0x86f7 */
            {8'h00}, /* 0x86f6 */
            {8'h00}, /* 0x86f5 */
            {8'h00}, /* 0x86f4 */
            {8'h00}, /* 0x86f3 */
            {8'h00}, /* 0x86f2 */
            {8'h00}, /* 0x86f1 */
            {8'h00}, /* 0x86f0 */
            {8'h00}, /* 0x86ef */
            {8'h00}, /* 0x86ee */
            {8'h00}, /* 0x86ed */
            {8'h00}, /* 0x86ec */
            {8'h00}, /* 0x86eb */
            {8'h00}, /* 0x86ea */
            {8'h00}, /* 0x86e9 */
            {8'h00}, /* 0x86e8 */
            {8'h00}, /* 0x86e7 */
            {8'h00}, /* 0x86e6 */
            {8'h00}, /* 0x86e5 */
            {8'h00}, /* 0x86e4 */
            {8'h00}, /* 0x86e3 */
            {8'h00}, /* 0x86e2 */
            {8'h00}, /* 0x86e1 */
            {8'h00}, /* 0x86e0 */
            {8'h00}, /* 0x86df */
            {8'h00}, /* 0x86de */
            {8'h00}, /* 0x86dd */
            {8'h00}, /* 0x86dc */
            {8'h00}, /* 0x86db */
            {8'h00}, /* 0x86da */
            {8'h00}, /* 0x86d9 */
            {8'h00}, /* 0x86d8 */
            {8'h00}, /* 0x86d7 */
            {8'h00}, /* 0x86d6 */
            {8'h00}, /* 0x86d5 */
            {8'h00}, /* 0x86d4 */
            {8'h00}, /* 0x86d3 */
            {8'h00}, /* 0x86d2 */
            {8'h00}, /* 0x86d1 */
            {8'h00}, /* 0x86d0 */
            {8'h00}, /* 0x86cf */
            {8'h00}, /* 0x86ce */
            {8'h00}, /* 0x86cd */
            {8'h00}, /* 0x86cc */
            {8'h00}, /* 0x86cb */
            {8'h00}, /* 0x86ca */
            {8'h00}, /* 0x86c9 */
            {8'h00}, /* 0x86c8 */
            {8'h00}, /* 0x86c7 */
            {8'h00}, /* 0x86c6 */
            {8'h00}, /* 0x86c5 */
            {8'h00}, /* 0x86c4 */
            {8'h00}, /* 0x86c3 */
            {8'h00}, /* 0x86c2 */
            {8'h00}, /* 0x86c1 */
            {8'h00}, /* 0x86c0 */
            {8'h00}, /* 0x86bf */
            {8'h00}, /* 0x86be */
            {8'h00}, /* 0x86bd */
            {8'h00}, /* 0x86bc */
            {8'h00}, /* 0x86bb */
            {8'h00}, /* 0x86ba */
            {8'h00}, /* 0x86b9 */
            {8'h00}, /* 0x86b8 */
            {8'h00}, /* 0x86b7 */
            {8'h00}, /* 0x86b6 */
            {8'h00}, /* 0x86b5 */
            {8'h00}, /* 0x86b4 */
            {8'h00}, /* 0x86b3 */
            {8'h00}, /* 0x86b2 */
            {8'h00}, /* 0x86b1 */
            {8'h00}, /* 0x86b0 */
            {8'h00}, /* 0x86af */
            {8'h00}, /* 0x86ae */
            {8'h00}, /* 0x86ad */
            {8'h00}, /* 0x86ac */
            {8'h00}, /* 0x86ab */
            {8'h00}, /* 0x86aa */
            {8'h00}, /* 0x86a9 */
            {8'h00}, /* 0x86a8 */
            {8'h00}, /* 0x86a7 */
            {8'h00}, /* 0x86a6 */
            {8'h00}, /* 0x86a5 */
            {8'h00}, /* 0x86a4 */
            {8'h00}, /* 0x86a3 */
            {8'h00}, /* 0x86a2 */
            {8'h00}, /* 0x86a1 */
            {8'h00}, /* 0x86a0 */
            {8'h00}, /* 0x869f */
            {8'h00}, /* 0x869e */
            {8'h00}, /* 0x869d */
            {8'h00}, /* 0x869c */
            {8'h00}, /* 0x869b */
            {8'h00}, /* 0x869a */
            {8'h00}, /* 0x8699 */
            {8'h00}, /* 0x8698 */
            {8'h00}, /* 0x8697 */
            {8'h00}, /* 0x8696 */
            {8'h00}, /* 0x8695 */
            {8'h00}, /* 0x8694 */
            {8'h00}, /* 0x8693 */
            {8'h00}, /* 0x8692 */
            {8'h00}, /* 0x8691 */
            {8'h00}, /* 0x8690 */
            {8'h00}, /* 0x868f */
            {8'h00}, /* 0x868e */
            {8'h00}, /* 0x868d */
            {8'h00}, /* 0x868c */
            {8'h00}, /* 0x868b */
            {8'h00}, /* 0x868a */
            {8'h00}, /* 0x8689 */
            {8'h00}, /* 0x8688 */
            {8'h00}, /* 0x8687 */
            {8'h00}, /* 0x8686 */
            {8'h00}, /* 0x8685 */
            {8'h00}, /* 0x8684 */
            {8'h00}, /* 0x8683 */
            {8'h00}, /* 0x8682 */
            {8'h00}, /* 0x8681 */
            {8'h00}, /* 0x8680 */
            {8'h00}, /* 0x867f */
            {8'h00}, /* 0x867e */
            {8'h00}, /* 0x867d */
            {8'h00}, /* 0x867c */
            {8'h00}, /* 0x867b */
            {8'h00}, /* 0x867a */
            {8'h00}, /* 0x8679 */
            {8'h00}, /* 0x8678 */
            {8'h00}, /* 0x8677 */
            {8'h00}, /* 0x8676 */
            {8'h00}, /* 0x8675 */
            {8'h00}, /* 0x8674 */
            {8'h00}, /* 0x8673 */
            {8'h00}, /* 0x8672 */
            {8'h00}, /* 0x8671 */
            {8'h00}, /* 0x8670 */
            {8'h00}, /* 0x866f */
            {8'h00}, /* 0x866e */
            {8'h00}, /* 0x866d */
            {8'h00}, /* 0x866c */
            {8'h00}, /* 0x866b */
            {8'h00}, /* 0x866a */
            {8'h00}, /* 0x8669 */
            {8'h00}, /* 0x8668 */
            {8'h00}, /* 0x8667 */
            {8'h00}, /* 0x8666 */
            {8'h00}, /* 0x8665 */
            {8'h00}, /* 0x8664 */
            {8'h00}, /* 0x8663 */
            {8'h00}, /* 0x8662 */
            {8'h00}, /* 0x8661 */
            {8'h00}, /* 0x8660 */
            {8'h00}, /* 0x865f */
            {8'h00}, /* 0x865e */
            {8'h00}, /* 0x865d */
            {8'h00}, /* 0x865c */
            {8'h00}, /* 0x865b */
            {8'h00}, /* 0x865a */
            {8'h00}, /* 0x8659 */
            {8'h00}, /* 0x8658 */
            {8'h00}, /* 0x8657 */
            {8'h00}, /* 0x8656 */
            {8'h00}, /* 0x8655 */
            {8'h00}, /* 0x8654 */
            {8'h00}, /* 0x8653 */
            {8'h00}, /* 0x8652 */
            {8'h00}, /* 0x8651 */
            {8'h00}, /* 0x8650 */
            {8'h00}, /* 0x864f */
            {8'h00}, /* 0x864e */
            {8'h00}, /* 0x864d */
            {8'h00}, /* 0x864c */
            {8'h00}, /* 0x864b */
            {8'h00}, /* 0x864a */
            {8'h00}, /* 0x8649 */
            {8'h00}, /* 0x8648 */
            {8'h00}, /* 0x8647 */
            {8'h00}, /* 0x8646 */
            {8'h00}, /* 0x8645 */
            {8'h00}, /* 0x8644 */
            {8'h00}, /* 0x8643 */
            {8'h00}, /* 0x8642 */
            {8'h00}, /* 0x8641 */
            {8'h00}, /* 0x8640 */
            {8'h00}, /* 0x863f */
            {8'h00}, /* 0x863e */
            {8'h00}, /* 0x863d */
            {8'h00}, /* 0x863c */
            {8'h00}, /* 0x863b */
            {8'h00}, /* 0x863a */
            {8'h00}, /* 0x8639 */
            {8'h00}, /* 0x8638 */
            {8'h00}, /* 0x8637 */
            {8'h00}, /* 0x8636 */
            {8'h00}, /* 0x8635 */
            {8'h00}, /* 0x8634 */
            {8'h00}, /* 0x8633 */
            {8'h00}, /* 0x8632 */
            {8'h00}, /* 0x8631 */
            {8'h00}, /* 0x8630 */
            {8'h00}, /* 0x862f */
            {8'h00}, /* 0x862e */
            {8'h00}, /* 0x862d */
            {8'h00}, /* 0x862c */
            {8'h00}, /* 0x862b */
            {8'h00}, /* 0x862a */
            {8'h00}, /* 0x8629 */
            {8'h00}, /* 0x8628 */
            {8'h00}, /* 0x8627 */
            {8'h00}, /* 0x8626 */
            {8'h00}, /* 0x8625 */
            {8'h00}, /* 0x8624 */
            {8'h00}, /* 0x8623 */
            {8'h00}, /* 0x8622 */
            {8'h00}, /* 0x8621 */
            {8'h00}, /* 0x8620 */
            {8'h00}, /* 0x861f */
            {8'h00}, /* 0x861e */
            {8'h00}, /* 0x861d */
            {8'h00}, /* 0x861c */
            {8'h00}, /* 0x861b */
            {8'h00}, /* 0x861a */
            {8'h00}, /* 0x8619 */
            {8'h00}, /* 0x8618 */
            {8'h00}, /* 0x8617 */
            {8'h00}, /* 0x8616 */
            {8'h00}, /* 0x8615 */
            {8'h00}, /* 0x8614 */
            {8'h00}, /* 0x8613 */
            {8'h00}, /* 0x8612 */
            {8'h00}, /* 0x8611 */
            {8'h00}, /* 0x8610 */
            {8'h00}, /* 0x860f */
            {8'h00}, /* 0x860e */
            {8'h00}, /* 0x860d */
            {8'h00}, /* 0x860c */
            {8'h00}, /* 0x860b */
            {8'h00}, /* 0x860a */
            {8'h00}, /* 0x8609 */
            {8'h00}, /* 0x8608 */
            {8'h00}, /* 0x8607 */
            {8'h00}, /* 0x8606 */
            {8'h00}, /* 0x8605 */
            {8'h00}, /* 0x8604 */
            {8'h00}, /* 0x8603 */
            {8'h00}, /* 0x8602 */
            {8'h00}, /* 0x8601 */
            {8'h00}, /* 0x8600 */
            {8'h00}, /* 0x85ff */
            {8'h00}, /* 0x85fe */
            {8'h00}, /* 0x85fd */
            {8'h00}, /* 0x85fc */
            {8'h00}, /* 0x85fb */
            {8'h00}, /* 0x85fa */
            {8'h00}, /* 0x85f9 */
            {8'h00}, /* 0x85f8 */
            {8'h00}, /* 0x85f7 */
            {8'h00}, /* 0x85f6 */
            {8'h00}, /* 0x85f5 */
            {8'h00}, /* 0x85f4 */
            {8'h00}, /* 0x85f3 */
            {8'h00}, /* 0x85f2 */
            {8'h00}, /* 0x85f1 */
            {8'h00}, /* 0x85f0 */
            {8'h00}, /* 0x85ef */
            {8'h00}, /* 0x85ee */
            {8'h00}, /* 0x85ed */
            {8'h00}, /* 0x85ec */
            {8'h00}, /* 0x85eb */
            {8'h00}, /* 0x85ea */
            {8'h00}, /* 0x85e9 */
            {8'h00}, /* 0x85e8 */
            {8'h00}, /* 0x85e7 */
            {8'h00}, /* 0x85e6 */
            {8'h00}, /* 0x85e5 */
            {8'h00}, /* 0x85e4 */
            {8'h00}, /* 0x85e3 */
            {8'h00}, /* 0x85e2 */
            {8'h00}, /* 0x85e1 */
            {8'h00}, /* 0x85e0 */
            {8'h00}, /* 0x85df */
            {8'h00}, /* 0x85de */
            {8'h00}, /* 0x85dd */
            {8'h00}, /* 0x85dc */
            {8'h00}, /* 0x85db */
            {8'h00}, /* 0x85da */
            {8'h00}, /* 0x85d9 */
            {8'h00}, /* 0x85d8 */
            {8'h00}, /* 0x85d7 */
            {8'h00}, /* 0x85d6 */
            {8'h00}, /* 0x85d5 */
            {8'h00}, /* 0x85d4 */
            {8'h00}, /* 0x85d3 */
            {8'h00}, /* 0x85d2 */
            {8'h00}, /* 0x85d1 */
            {8'h00}, /* 0x85d0 */
            {8'h00}, /* 0x85cf */
            {8'h00}, /* 0x85ce */
            {8'h00}, /* 0x85cd */
            {8'h00}, /* 0x85cc */
            {8'h00}, /* 0x85cb */
            {8'h00}, /* 0x85ca */
            {8'h00}, /* 0x85c9 */
            {8'h00}, /* 0x85c8 */
            {8'h00}, /* 0x85c7 */
            {8'h00}, /* 0x85c6 */
            {8'h00}, /* 0x85c5 */
            {8'h00}, /* 0x85c4 */
            {8'h00}, /* 0x85c3 */
            {8'h00}, /* 0x85c2 */
            {8'h00}, /* 0x85c1 */
            {8'h00}, /* 0x85c0 */
            {8'h00}, /* 0x85bf */
            {8'h00}, /* 0x85be */
            {8'h00}, /* 0x85bd */
            {8'h00}, /* 0x85bc */
            {8'h00}, /* 0x85bb */
            {8'h00}, /* 0x85ba */
            {8'h00}, /* 0x85b9 */
            {8'h00}, /* 0x85b8 */
            {8'h00}, /* 0x85b7 */
            {8'h00}, /* 0x85b6 */
            {8'h00}, /* 0x85b5 */
            {8'h00}, /* 0x85b4 */
            {8'h00}, /* 0x85b3 */
            {8'h00}, /* 0x85b2 */
            {8'h00}, /* 0x85b1 */
            {8'h00}, /* 0x85b0 */
            {8'h00}, /* 0x85af */
            {8'h00}, /* 0x85ae */
            {8'h00}, /* 0x85ad */
            {8'h00}, /* 0x85ac */
            {8'h00}, /* 0x85ab */
            {8'h00}, /* 0x85aa */
            {8'h00}, /* 0x85a9 */
            {8'h00}, /* 0x85a8 */
            {8'h00}, /* 0x85a7 */
            {8'h00}, /* 0x85a6 */
            {8'h00}, /* 0x85a5 */
            {8'h00}, /* 0x85a4 */
            {8'h00}, /* 0x85a3 */
            {8'h00}, /* 0x85a2 */
            {8'h00}, /* 0x85a1 */
            {8'h00}, /* 0x85a0 */
            {8'h00}, /* 0x859f */
            {8'h00}, /* 0x859e */
            {8'h00}, /* 0x859d */
            {8'h00}, /* 0x859c */
            {8'h00}, /* 0x859b */
            {8'h00}, /* 0x859a */
            {8'h00}, /* 0x8599 */
            {8'h00}, /* 0x8598 */
            {8'h00}, /* 0x8597 */
            {8'h00}, /* 0x8596 */
            {8'h00}, /* 0x8595 */
            {8'h00}, /* 0x8594 */
            {8'h00}, /* 0x8593 */
            {8'h00}, /* 0x8592 */
            {8'h00}, /* 0x8591 */
            {8'h00}, /* 0x8590 */
            {8'h00}, /* 0x858f */
            {8'h00}, /* 0x858e */
            {8'h00}, /* 0x858d */
            {8'h00}, /* 0x858c */
            {8'h00}, /* 0x858b */
            {8'h00}, /* 0x858a */
            {8'h00}, /* 0x8589 */
            {8'h00}, /* 0x8588 */
            {8'h00}, /* 0x8587 */
            {8'h00}, /* 0x8586 */
            {8'h00}, /* 0x8585 */
            {8'h00}, /* 0x8584 */
            {8'h00}, /* 0x8583 */
            {8'h00}, /* 0x8582 */
            {8'h00}, /* 0x8581 */
            {8'h00}, /* 0x8580 */
            {8'h00}, /* 0x857f */
            {8'h00}, /* 0x857e */
            {8'h00}, /* 0x857d */
            {8'h00}, /* 0x857c */
            {8'h00}, /* 0x857b */
            {8'h00}, /* 0x857a */
            {8'h00}, /* 0x8579 */
            {8'h00}, /* 0x8578 */
            {8'h00}, /* 0x8577 */
            {8'h00}, /* 0x8576 */
            {8'h00}, /* 0x8575 */
            {8'h00}, /* 0x8574 */
            {8'h00}, /* 0x8573 */
            {8'h00}, /* 0x8572 */
            {8'h00}, /* 0x8571 */
            {8'h00}, /* 0x8570 */
            {8'h00}, /* 0x856f */
            {8'h00}, /* 0x856e */
            {8'h00}, /* 0x856d */
            {8'h00}, /* 0x856c */
            {8'h00}, /* 0x856b */
            {8'h00}, /* 0x856a */
            {8'h00}, /* 0x8569 */
            {8'h00}, /* 0x8568 */
            {8'h00}, /* 0x8567 */
            {8'h00}, /* 0x8566 */
            {8'h00}, /* 0x8565 */
            {8'h00}, /* 0x8564 */
            {8'h00}, /* 0x8563 */
            {8'h00}, /* 0x8562 */
            {8'h00}, /* 0x8561 */
            {8'h00}, /* 0x8560 */
            {8'h00}, /* 0x855f */
            {8'h00}, /* 0x855e */
            {8'h00}, /* 0x855d */
            {8'h00}, /* 0x855c */
            {8'h00}, /* 0x855b */
            {8'h00}, /* 0x855a */
            {8'h00}, /* 0x8559 */
            {8'h00}, /* 0x8558 */
            {8'h00}, /* 0x8557 */
            {8'h00}, /* 0x8556 */
            {8'h00}, /* 0x8555 */
            {8'h00}, /* 0x8554 */
            {8'h00}, /* 0x8553 */
            {8'h00}, /* 0x8552 */
            {8'h00}, /* 0x8551 */
            {8'h00}, /* 0x8550 */
            {8'h00}, /* 0x854f */
            {8'h00}, /* 0x854e */
            {8'h00}, /* 0x854d */
            {8'h00}, /* 0x854c */
            {8'h00}, /* 0x854b */
            {8'h00}, /* 0x854a */
            {8'h00}, /* 0x8549 */
            {8'h00}, /* 0x8548 */
            {8'h00}, /* 0x8547 */
            {8'h00}, /* 0x8546 */
            {8'h00}, /* 0x8545 */
            {8'h00}, /* 0x8544 */
            {8'h00}, /* 0x8543 */
            {8'h00}, /* 0x8542 */
            {8'h00}, /* 0x8541 */
            {8'h00}, /* 0x8540 */
            {8'h00}, /* 0x853f */
            {8'h00}, /* 0x853e */
            {8'h00}, /* 0x853d */
            {8'h00}, /* 0x853c */
            {8'h00}, /* 0x853b */
            {8'h00}, /* 0x853a */
            {8'h00}, /* 0x8539 */
            {8'h00}, /* 0x8538 */
            {8'h00}, /* 0x8537 */
            {8'h00}, /* 0x8536 */
            {8'h00}, /* 0x8535 */
            {8'h00}, /* 0x8534 */
            {8'h00}, /* 0x8533 */
            {8'h00}, /* 0x8532 */
            {8'h00}, /* 0x8531 */
            {8'h00}, /* 0x8530 */
            {8'h00}, /* 0x852f */
            {8'h00}, /* 0x852e */
            {8'h00}, /* 0x852d */
            {8'h00}, /* 0x852c */
            {8'h00}, /* 0x852b */
            {8'h00}, /* 0x852a */
            {8'h00}, /* 0x8529 */
            {8'h00}, /* 0x8528 */
            {8'h00}, /* 0x8527 */
            {8'h00}, /* 0x8526 */
            {8'h00}, /* 0x8525 */
            {8'h00}, /* 0x8524 */
            {8'h00}, /* 0x8523 */
            {8'h00}, /* 0x8522 */
            {8'h00}, /* 0x8521 */
            {8'h00}, /* 0x8520 */
            {8'h00}, /* 0x851f */
            {8'h00}, /* 0x851e */
            {8'h00}, /* 0x851d */
            {8'h00}, /* 0x851c */
            {8'h00}, /* 0x851b */
            {8'h00}, /* 0x851a */
            {8'h00}, /* 0x8519 */
            {8'h00}, /* 0x8518 */
            {8'h00}, /* 0x8517 */
            {8'h00}, /* 0x8516 */
            {8'h00}, /* 0x8515 */
            {8'h00}, /* 0x8514 */
            {8'h00}, /* 0x8513 */
            {8'h00}, /* 0x8512 */
            {8'h00}, /* 0x8511 */
            {8'h00}, /* 0x8510 */
            {8'h00}, /* 0x850f */
            {8'h00}, /* 0x850e */
            {8'h00}, /* 0x850d */
            {8'h00}, /* 0x850c */
            {8'h00}, /* 0x850b */
            {8'h00}, /* 0x850a */
            {8'h00}, /* 0x8509 */
            {8'h00}, /* 0x8508 */
            {8'h00}, /* 0x8507 */
            {8'h00}, /* 0x8506 */
            {8'h00}, /* 0x8505 */
            {8'h00}, /* 0x8504 */
            {8'h00}, /* 0x8503 */
            {8'h00}, /* 0x8502 */
            {8'h00}, /* 0x8501 */
            {8'h00}, /* 0x8500 */
            {8'h00}, /* 0x84ff */
            {8'h00}, /* 0x84fe */
            {8'h00}, /* 0x84fd */
            {8'h00}, /* 0x84fc */
            {8'h00}, /* 0x84fb */
            {8'h00}, /* 0x84fa */
            {8'h00}, /* 0x84f9 */
            {8'h00}, /* 0x84f8 */
            {8'h00}, /* 0x84f7 */
            {8'h00}, /* 0x84f6 */
            {8'h00}, /* 0x84f5 */
            {8'h00}, /* 0x84f4 */
            {8'h00}, /* 0x84f3 */
            {8'h00}, /* 0x84f2 */
            {8'h00}, /* 0x84f1 */
            {8'h00}, /* 0x84f0 */
            {8'h00}, /* 0x84ef */
            {8'h00}, /* 0x84ee */
            {8'h00}, /* 0x84ed */
            {8'h00}, /* 0x84ec */
            {8'h00}, /* 0x84eb */
            {8'h00}, /* 0x84ea */
            {8'h00}, /* 0x84e9 */
            {8'h00}, /* 0x84e8 */
            {8'h00}, /* 0x84e7 */
            {8'h00}, /* 0x84e6 */
            {8'h00}, /* 0x84e5 */
            {8'h00}, /* 0x84e4 */
            {8'h00}, /* 0x84e3 */
            {8'h00}, /* 0x84e2 */
            {8'h00}, /* 0x84e1 */
            {8'h00}, /* 0x84e0 */
            {8'h00}, /* 0x84df */
            {8'h00}, /* 0x84de */
            {8'h00}, /* 0x84dd */
            {8'h00}, /* 0x84dc */
            {8'h00}, /* 0x84db */
            {8'h00}, /* 0x84da */
            {8'h00}, /* 0x84d9 */
            {8'h00}, /* 0x84d8 */
            {8'h00}, /* 0x84d7 */
            {8'h00}, /* 0x84d6 */
            {8'h00}, /* 0x84d5 */
            {8'h00}, /* 0x84d4 */
            {8'h00}, /* 0x84d3 */
            {8'h00}, /* 0x84d2 */
            {8'h00}, /* 0x84d1 */
            {8'h00}, /* 0x84d0 */
            {8'h00}, /* 0x84cf */
            {8'h00}, /* 0x84ce */
            {8'h00}, /* 0x84cd */
            {8'h00}, /* 0x84cc */
            {8'h00}, /* 0x84cb */
            {8'h00}, /* 0x84ca */
            {8'h00}, /* 0x84c9 */
            {8'h00}, /* 0x84c8 */
            {8'h00}, /* 0x84c7 */
            {8'h00}, /* 0x84c6 */
            {8'h00}, /* 0x84c5 */
            {8'h00}, /* 0x84c4 */
            {8'h00}, /* 0x84c3 */
            {8'h00}, /* 0x84c2 */
            {8'h00}, /* 0x84c1 */
            {8'h00}, /* 0x84c0 */
            {8'h00}, /* 0x84bf */
            {8'h00}, /* 0x84be */
            {8'h00}, /* 0x84bd */
            {8'h00}, /* 0x84bc */
            {8'h00}, /* 0x84bb */
            {8'h00}, /* 0x84ba */
            {8'h00}, /* 0x84b9 */
            {8'h00}, /* 0x84b8 */
            {8'h00}, /* 0x84b7 */
            {8'h00}, /* 0x84b6 */
            {8'h00}, /* 0x84b5 */
            {8'h00}, /* 0x84b4 */
            {8'h00}, /* 0x84b3 */
            {8'h00}, /* 0x84b2 */
            {8'h00}, /* 0x84b1 */
            {8'h00}, /* 0x84b0 */
            {8'h00}, /* 0x84af */
            {8'h00}, /* 0x84ae */
            {8'h00}, /* 0x84ad */
            {8'h00}, /* 0x84ac */
            {8'h00}, /* 0x84ab */
            {8'h00}, /* 0x84aa */
            {8'h00}, /* 0x84a9 */
            {8'h00}, /* 0x84a8 */
            {8'h00}, /* 0x84a7 */
            {8'h00}, /* 0x84a6 */
            {8'h00}, /* 0x84a5 */
            {8'h00}, /* 0x84a4 */
            {8'h00}, /* 0x84a3 */
            {8'h00}, /* 0x84a2 */
            {8'h00}, /* 0x84a1 */
            {8'h00}, /* 0x84a0 */
            {8'h00}, /* 0x849f */
            {8'h00}, /* 0x849e */
            {8'h00}, /* 0x849d */
            {8'h00}, /* 0x849c */
            {8'h00}, /* 0x849b */
            {8'h00}, /* 0x849a */
            {8'h00}, /* 0x8499 */
            {8'h00}, /* 0x8498 */
            {8'h00}, /* 0x8497 */
            {8'h00}, /* 0x8496 */
            {8'h00}, /* 0x8495 */
            {8'h00}, /* 0x8494 */
            {8'h00}, /* 0x8493 */
            {8'h00}, /* 0x8492 */
            {8'h00}, /* 0x8491 */
            {8'h00}, /* 0x8490 */
            {8'h00}, /* 0x848f */
            {8'h00}, /* 0x848e */
            {8'h00}, /* 0x848d */
            {8'h00}, /* 0x848c */
            {8'h00}, /* 0x848b */
            {8'h00}, /* 0x848a */
            {8'h00}, /* 0x8489 */
            {8'h00}, /* 0x8488 */
            {8'h00}, /* 0x8487 */
            {8'h00}, /* 0x8486 */
            {8'h00}, /* 0x8485 */
            {8'h00}, /* 0x8484 */
            {8'h00}, /* 0x8483 */
            {8'h00}, /* 0x8482 */
            {8'h00}, /* 0x8481 */
            {8'h00}, /* 0x8480 */
            {8'h00}, /* 0x847f */
            {8'h00}, /* 0x847e */
            {8'h00}, /* 0x847d */
            {8'h00}, /* 0x847c */
            {8'h00}, /* 0x847b */
            {8'h00}, /* 0x847a */
            {8'h00}, /* 0x8479 */
            {8'h00}, /* 0x8478 */
            {8'h00}, /* 0x8477 */
            {8'h00}, /* 0x8476 */
            {8'h00}, /* 0x8475 */
            {8'h00}, /* 0x8474 */
            {8'h00}, /* 0x8473 */
            {8'h00}, /* 0x8472 */
            {8'h00}, /* 0x8471 */
            {8'h00}, /* 0x8470 */
            {8'h00}, /* 0x846f */
            {8'h00}, /* 0x846e */
            {8'h00}, /* 0x846d */
            {8'h00}, /* 0x846c */
            {8'h00}, /* 0x846b */
            {8'h00}, /* 0x846a */
            {8'h00}, /* 0x8469 */
            {8'h00}, /* 0x8468 */
            {8'h00}, /* 0x8467 */
            {8'h00}, /* 0x8466 */
            {8'h00}, /* 0x8465 */
            {8'h00}, /* 0x8464 */
            {8'h00}, /* 0x8463 */
            {8'h00}, /* 0x8462 */
            {8'h00}, /* 0x8461 */
            {8'h00}, /* 0x8460 */
            {8'h00}, /* 0x845f */
            {8'h00}, /* 0x845e */
            {8'h00}, /* 0x845d */
            {8'h00}, /* 0x845c */
            {8'h00}, /* 0x845b */
            {8'h00}, /* 0x845a */
            {8'h00}, /* 0x8459 */
            {8'h00}, /* 0x8458 */
            {8'h00}, /* 0x8457 */
            {8'h00}, /* 0x8456 */
            {8'h00}, /* 0x8455 */
            {8'h00}, /* 0x8454 */
            {8'h00}, /* 0x8453 */
            {8'h00}, /* 0x8452 */
            {8'h00}, /* 0x8451 */
            {8'h00}, /* 0x8450 */
            {8'h00}, /* 0x844f */
            {8'h00}, /* 0x844e */
            {8'h00}, /* 0x844d */
            {8'h00}, /* 0x844c */
            {8'h00}, /* 0x844b */
            {8'h00}, /* 0x844a */
            {8'h00}, /* 0x8449 */
            {8'h00}, /* 0x8448 */
            {8'h00}, /* 0x8447 */
            {8'h00}, /* 0x8446 */
            {8'h00}, /* 0x8445 */
            {8'h00}, /* 0x8444 */
            {8'h00}, /* 0x8443 */
            {8'h00}, /* 0x8442 */
            {8'h00}, /* 0x8441 */
            {8'h00}, /* 0x8440 */
            {8'h00}, /* 0x843f */
            {8'h00}, /* 0x843e */
            {8'h00}, /* 0x843d */
            {8'h00}, /* 0x843c */
            {8'h00}, /* 0x843b */
            {8'h00}, /* 0x843a */
            {8'h00}, /* 0x8439 */
            {8'h00}, /* 0x8438 */
            {8'h00}, /* 0x8437 */
            {8'h00}, /* 0x8436 */
            {8'h00}, /* 0x8435 */
            {8'h00}, /* 0x8434 */
            {8'h00}, /* 0x8433 */
            {8'h00}, /* 0x8432 */
            {8'h00}, /* 0x8431 */
            {8'h00}, /* 0x8430 */
            {8'h00}, /* 0x842f */
            {8'h00}, /* 0x842e */
            {8'h00}, /* 0x842d */
            {8'h00}, /* 0x842c */
            {8'h00}, /* 0x842b */
            {8'h00}, /* 0x842a */
            {8'h00}, /* 0x8429 */
            {8'h00}, /* 0x8428 */
            {8'h00}, /* 0x8427 */
            {8'h00}, /* 0x8426 */
            {8'h00}, /* 0x8425 */
            {8'h00}, /* 0x8424 */
            {8'h00}, /* 0x8423 */
            {8'h00}, /* 0x8422 */
            {8'h00}, /* 0x8421 */
            {8'h00}, /* 0x8420 */
            {8'h00}, /* 0x841f */
            {8'h00}, /* 0x841e */
            {8'h00}, /* 0x841d */
            {8'h00}, /* 0x841c */
            {8'h00}, /* 0x841b */
            {8'h00}, /* 0x841a */
            {8'h00}, /* 0x8419 */
            {8'h00}, /* 0x8418 */
            {8'h00}, /* 0x8417 */
            {8'h00}, /* 0x8416 */
            {8'h00}, /* 0x8415 */
            {8'h00}, /* 0x8414 */
            {8'h00}, /* 0x8413 */
            {8'h00}, /* 0x8412 */
            {8'h00}, /* 0x8411 */
            {8'h00}, /* 0x8410 */
            {8'h00}, /* 0x840f */
            {8'h00}, /* 0x840e */
            {8'h00}, /* 0x840d */
            {8'h00}, /* 0x840c */
            {8'h00}, /* 0x840b */
            {8'h00}, /* 0x840a */
            {8'h00}, /* 0x8409 */
            {8'h00}, /* 0x8408 */
            {8'h00}, /* 0x8407 */
            {8'h00}, /* 0x8406 */
            {8'h00}, /* 0x8405 */
            {8'h00}, /* 0x8404 */
            {8'h00}, /* 0x8403 */
            {8'h00}, /* 0x8402 */
            {8'h00}, /* 0x8401 */
            {8'h00}, /* 0x8400 */
            {8'h00}, /* 0x83ff */
            {8'h00}, /* 0x83fe */
            {8'h00}, /* 0x83fd */
            {8'h00}, /* 0x83fc */
            {8'h00}, /* 0x83fb */
            {8'h00}, /* 0x83fa */
            {8'h00}, /* 0x83f9 */
            {8'h00}, /* 0x83f8 */
            {8'h00}, /* 0x83f7 */
            {8'h00}, /* 0x83f6 */
            {8'h00}, /* 0x83f5 */
            {8'h00}, /* 0x83f4 */
            {8'h00}, /* 0x83f3 */
            {8'h00}, /* 0x83f2 */
            {8'h00}, /* 0x83f1 */
            {8'h00}, /* 0x83f0 */
            {8'h00}, /* 0x83ef */
            {8'h00}, /* 0x83ee */
            {8'h00}, /* 0x83ed */
            {8'h00}, /* 0x83ec */
            {8'h00}, /* 0x83eb */
            {8'h00}, /* 0x83ea */
            {8'h00}, /* 0x83e9 */
            {8'h00}, /* 0x83e8 */
            {8'h00}, /* 0x83e7 */
            {8'h00}, /* 0x83e6 */
            {8'h00}, /* 0x83e5 */
            {8'h00}, /* 0x83e4 */
            {8'h00}, /* 0x83e3 */
            {8'h00}, /* 0x83e2 */
            {8'h00}, /* 0x83e1 */
            {8'h00}, /* 0x83e0 */
            {8'h00}, /* 0x83df */
            {8'h00}, /* 0x83de */
            {8'h00}, /* 0x83dd */
            {8'h00}, /* 0x83dc */
            {8'h00}, /* 0x83db */
            {8'h00}, /* 0x83da */
            {8'h00}, /* 0x83d9 */
            {8'h00}, /* 0x83d8 */
            {8'h00}, /* 0x83d7 */
            {8'h00}, /* 0x83d6 */
            {8'h00}, /* 0x83d5 */
            {8'h00}, /* 0x83d4 */
            {8'h00}, /* 0x83d3 */
            {8'h00}, /* 0x83d2 */
            {8'h00}, /* 0x83d1 */
            {8'h00}, /* 0x83d0 */
            {8'h00}, /* 0x83cf */
            {8'h00}, /* 0x83ce */
            {8'h00}, /* 0x83cd */
            {8'h00}, /* 0x83cc */
            {8'h00}, /* 0x83cb */
            {8'h00}, /* 0x83ca */
            {8'h00}, /* 0x83c9 */
            {8'h00}, /* 0x83c8 */
            {8'h00}, /* 0x83c7 */
            {8'h00}, /* 0x83c6 */
            {8'h00}, /* 0x83c5 */
            {8'h00}, /* 0x83c4 */
            {8'h00}, /* 0x83c3 */
            {8'h00}, /* 0x83c2 */
            {8'h00}, /* 0x83c1 */
            {8'h00}, /* 0x83c0 */
            {8'h00}, /* 0x83bf */
            {8'h00}, /* 0x83be */
            {8'h00}, /* 0x83bd */
            {8'h00}, /* 0x83bc */
            {8'h00}, /* 0x83bb */
            {8'h00}, /* 0x83ba */
            {8'h00}, /* 0x83b9 */
            {8'h00}, /* 0x83b8 */
            {8'h00}, /* 0x83b7 */
            {8'h00}, /* 0x83b6 */
            {8'h00}, /* 0x83b5 */
            {8'h00}, /* 0x83b4 */
            {8'h00}, /* 0x83b3 */
            {8'h00}, /* 0x83b2 */
            {8'h00}, /* 0x83b1 */
            {8'h00}, /* 0x83b0 */
            {8'h00}, /* 0x83af */
            {8'h00}, /* 0x83ae */
            {8'h00}, /* 0x83ad */
            {8'h00}, /* 0x83ac */
            {8'h00}, /* 0x83ab */
            {8'h00}, /* 0x83aa */
            {8'h00}, /* 0x83a9 */
            {8'h00}, /* 0x83a8 */
            {8'h00}, /* 0x83a7 */
            {8'h00}, /* 0x83a6 */
            {8'h00}, /* 0x83a5 */
            {8'h00}, /* 0x83a4 */
            {8'h00}, /* 0x83a3 */
            {8'h00}, /* 0x83a2 */
            {8'h00}, /* 0x83a1 */
            {8'h00}, /* 0x83a0 */
            {8'h00}, /* 0x839f */
            {8'h00}, /* 0x839e */
            {8'h00}, /* 0x839d */
            {8'h00}, /* 0x839c */
            {8'h00}, /* 0x839b */
            {8'h00}, /* 0x839a */
            {8'h00}, /* 0x8399 */
            {8'h00}, /* 0x8398 */
            {8'h00}, /* 0x8397 */
            {8'h00}, /* 0x8396 */
            {8'h00}, /* 0x8395 */
            {8'h00}, /* 0x8394 */
            {8'h00}, /* 0x8393 */
            {8'h00}, /* 0x8392 */
            {8'h00}, /* 0x8391 */
            {8'h00}, /* 0x8390 */
            {8'h00}, /* 0x838f */
            {8'h00}, /* 0x838e */
            {8'h00}, /* 0x838d */
            {8'h00}, /* 0x838c */
            {8'h00}, /* 0x838b */
            {8'h00}, /* 0x838a */
            {8'h00}, /* 0x8389 */
            {8'h00}, /* 0x8388 */
            {8'h00}, /* 0x8387 */
            {8'h00}, /* 0x8386 */
            {8'h00}, /* 0x8385 */
            {8'h00}, /* 0x8384 */
            {8'h00}, /* 0x8383 */
            {8'h00}, /* 0x8382 */
            {8'h00}, /* 0x8381 */
            {8'h00}, /* 0x8380 */
            {8'h00}, /* 0x837f */
            {8'h00}, /* 0x837e */
            {8'h00}, /* 0x837d */
            {8'h00}, /* 0x837c */
            {8'h00}, /* 0x837b */
            {8'h00}, /* 0x837a */
            {8'h00}, /* 0x8379 */
            {8'h00}, /* 0x8378 */
            {8'h00}, /* 0x8377 */
            {8'h00}, /* 0x8376 */
            {8'h00}, /* 0x8375 */
            {8'h00}, /* 0x8374 */
            {8'h00}, /* 0x8373 */
            {8'h00}, /* 0x8372 */
            {8'h00}, /* 0x8371 */
            {8'h00}, /* 0x8370 */
            {8'h00}, /* 0x836f */
            {8'h00}, /* 0x836e */
            {8'h00}, /* 0x836d */
            {8'h00}, /* 0x836c */
            {8'h00}, /* 0x836b */
            {8'h00}, /* 0x836a */
            {8'h00}, /* 0x8369 */
            {8'h00}, /* 0x8368 */
            {8'h00}, /* 0x8367 */
            {8'h00}, /* 0x8366 */
            {8'h00}, /* 0x8365 */
            {8'h00}, /* 0x8364 */
            {8'h00}, /* 0x8363 */
            {8'h00}, /* 0x8362 */
            {8'h00}, /* 0x8361 */
            {8'h00}, /* 0x8360 */
            {8'h00}, /* 0x835f */
            {8'h00}, /* 0x835e */
            {8'h00}, /* 0x835d */
            {8'h00}, /* 0x835c */
            {8'h00}, /* 0x835b */
            {8'h00}, /* 0x835a */
            {8'h00}, /* 0x8359 */
            {8'h00}, /* 0x8358 */
            {8'h00}, /* 0x8357 */
            {8'h00}, /* 0x8356 */
            {8'h00}, /* 0x8355 */
            {8'h00}, /* 0x8354 */
            {8'h00}, /* 0x8353 */
            {8'h00}, /* 0x8352 */
            {8'h00}, /* 0x8351 */
            {8'h00}, /* 0x8350 */
            {8'h00}, /* 0x834f */
            {8'h00}, /* 0x834e */
            {8'h00}, /* 0x834d */
            {8'h00}, /* 0x834c */
            {8'h00}, /* 0x834b */
            {8'h00}, /* 0x834a */
            {8'h00}, /* 0x8349 */
            {8'h00}, /* 0x8348 */
            {8'h00}, /* 0x8347 */
            {8'h00}, /* 0x8346 */
            {8'h00}, /* 0x8345 */
            {8'h00}, /* 0x8344 */
            {8'h00}, /* 0x8343 */
            {8'h00}, /* 0x8342 */
            {8'h00}, /* 0x8341 */
            {8'h00}, /* 0x8340 */
            {8'h00}, /* 0x833f */
            {8'h00}, /* 0x833e */
            {8'h00}, /* 0x833d */
            {8'h00}, /* 0x833c */
            {8'h00}, /* 0x833b */
            {8'h00}, /* 0x833a */
            {8'h00}, /* 0x8339 */
            {8'h00}, /* 0x8338 */
            {8'h00}, /* 0x8337 */
            {8'h00}, /* 0x8336 */
            {8'h00}, /* 0x8335 */
            {8'h00}, /* 0x8334 */
            {8'h00}, /* 0x8333 */
            {8'h00}, /* 0x8332 */
            {8'h00}, /* 0x8331 */
            {8'h00}, /* 0x8330 */
            {8'h00}, /* 0x832f */
            {8'h00}, /* 0x832e */
            {8'h00}, /* 0x832d */
            {8'h00}, /* 0x832c */
            {8'h00}, /* 0x832b */
            {8'h00}, /* 0x832a */
            {8'h00}, /* 0x8329 */
            {8'h00}, /* 0x8328 */
            {8'h00}, /* 0x8327 */
            {8'h00}, /* 0x8326 */
            {8'h00}, /* 0x8325 */
            {8'h00}, /* 0x8324 */
            {8'h00}, /* 0x8323 */
            {8'h00}, /* 0x8322 */
            {8'h00}, /* 0x8321 */
            {8'h00}, /* 0x8320 */
            {8'h00}, /* 0x831f */
            {8'h00}, /* 0x831e */
            {8'h00}, /* 0x831d */
            {8'h00}, /* 0x831c */
            {8'h00}, /* 0x831b */
            {8'h00}, /* 0x831a */
            {8'h00}, /* 0x8319 */
            {8'h00}, /* 0x8318 */
            {8'h00}, /* 0x8317 */
            {8'h00}, /* 0x8316 */
            {8'h00}, /* 0x8315 */
            {8'h00}, /* 0x8314 */
            {8'h00}, /* 0x8313 */
            {8'h00}, /* 0x8312 */
            {8'h00}, /* 0x8311 */
            {8'h00}, /* 0x8310 */
            {8'h00}, /* 0x830f */
            {8'h00}, /* 0x830e */
            {8'h00}, /* 0x830d */
            {8'h00}, /* 0x830c */
            {8'h00}, /* 0x830b */
            {8'h00}, /* 0x830a */
            {8'h00}, /* 0x8309 */
            {8'h00}, /* 0x8308 */
            {8'h00}, /* 0x8307 */
            {8'h00}, /* 0x8306 */
            {8'h00}, /* 0x8305 */
            {8'h00}, /* 0x8304 */
            {8'h00}, /* 0x8303 */
            {8'h00}, /* 0x8302 */
            {8'h00}, /* 0x8301 */
            {8'h00}, /* 0x8300 */
            {8'h00}, /* 0x82ff */
            {8'h00}, /* 0x82fe */
            {8'h00}, /* 0x82fd */
            {8'h00}, /* 0x82fc */
            {8'h00}, /* 0x82fb */
            {8'h00}, /* 0x82fa */
            {8'h00}, /* 0x82f9 */
            {8'h00}, /* 0x82f8 */
            {8'h00}, /* 0x82f7 */
            {8'h00}, /* 0x82f6 */
            {8'h00}, /* 0x82f5 */
            {8'h00}, /* 0x82f4 */
            {8'h00}, /* 0x82f3 */
            {8'h00}, /* 0x82f2 */
            {8'h00}, /* 0x82f1 */
            {8'h00}, /* 0x82f0 */
            {8'h00}, /* 0x82ef */
            {8'h00}, /* 0x82ee */
            {8'h00}, /* 0x82ed */
            {8'h00}, /* 0x82ec */
            {8'h00}, /* 0x82eb */
            {8'h00}, /* 0x82ea */
            {8'h00}, /* 0x82e9 */
            {8'h00}, /* 0x82e8 */
            {8'h00}, /* 0x82e7 */
            {8'h00}, /* 0x82e6 */
            {8'h00}, /* 0x82e5 */
            {8'h00}, /* 0x82e4 */
            {8'h00}, /* 0x82e3 */
            {8'h00}, /* 0x82e2 */
            {8'h00}, /* 0x82e1 */
            {8'h00}, /* 0x82e0 */
            {8'h00}, /* 0x82df */
            {8'h00}, /* 0x82de */
            {8'h00}, /* 0x82dd */
            {8'h00}, /* 0x82dc */
            {8'h00}, /* 0x82db */
            {8'h00}, /* 0x82da */
            {8'h00}, /* 0x82d9 */
            {8'h00}, /* 0x82d8 */
            {8'h00}, /* 0x82d7 */
            {8'h00}, /* 0x82d6 */
            {8'h00}, /* 0x82d5 */
            {8'h00}, /* 0x82d4 */
            {8'h00}, /* 0x82d3 */
            {8'h00}, /* 0x82d2 */
            {8'h00}, /* 0x82d1 */
            {8'h00}, /* 0x82d0 */
            {8'h00}, /* 0x82cf */
            {8'h00}, /* 0x82ce */
            {8'h00}, /* 0x82cd */
            {8'h00}, /* 0x82cc */
            {8'h00}, /* 0x82cb */
            {8'h00}, /* 0x82ca */
            {8'h00}, /* 0x82c9 */
            {8'h00}, /* 0x82c8 */
            {8'h00}, /* 0x82c7 */
            {8'h00}, /* 0x82c6 */
            {8'h00}, /* 0x82c5 */
            {8'h00}, /* 0x82c4 */
            {8'h00}, /* 0x82c3 */
            {8'h00}, /* 0x82c2 */
            {8'h00}, /* 0x82c1 */
            {8'h00}, /* 0x82c0 */
            {8'h00}, /* 0x82bf */
            {8'h00}, /* 0x82be */
            {8'h00}, /* 0x82bd */
            {8'h00}, /* 0x82bc */
            {8'h00}, /* 0x82bb */
            {8'h00}, /* 0x82ba */
            {8'h00}, /* 0x82b9 */
            {8'h00}, /* 0x82b8 */
            {8'h00}, /* 0x82b7 */
            {8'h00}, /* 0x82b6 */
            {8'h00}, /* 0x82b5 */
            {8'h00}, /* 0x82b4 */
            {8'h00}, /* 0x82b3 */
            {8'h00}, /* 0x82b2 */
            {8'h00}, /* 0x82b1 */
            {8'h00}, /* 0x82b0 */
            {8'h00}, /* 0x82af */
            {8'h00}, /* 0x82ae */
            {8'h00}, /* 0x82ad */
            {8'h00}, /* 0x82ac */
            {8'h00}, /* 0x82ab */
            {8'h00}, /* 0x82aa */
            {8'h00}, /* 0x82a9 */
            {8'h00}, /* 0x82a8 */
            {8'h00}, /* 0x82a7 */
            {8'h00}, /* 0x82a6 */
            {8'h00}, /* 0x82a5 */
            {8'h00}, /* 0x82a4 */
            {8'h00}, /* 0x82a3 */
            {8'h00}, /* 0x82a2 */
            {8'h00}, /* 0x82a1 */
            {8'h00}, /* 0x82a0 */
            {8'h00}, /* 0x829f */
            {8'h00}, /* 0x829e */
            {8'h00}, /* 0x829d */
            {8'h00}, /* 0x829c */
            {8'h00}, /* 0x829b */
            {8'h00}, /* 0x829a */
            {8'h00}, /* 0x8299 */
            {8'h00}, /* 0x8298 */
            {8'h00}, /* 0x8297 */
            {8'h00}, /* 0x8296 */
            {8'h00}, /* 0x8295 */
            {8'h00}, /* 0x8294 */
            {8'h00}, /* 0x8293 */
            {8'h00}, /* 0x8292 */
            {8'h00}, /* 0x8291 */
            {8'h00}, /* 0x8290 */
            {8'h00}, /* 0x828f */
            {8'h00}, /* 0x828e */
            {8'h00}, /* 0x828d */
            {8'h00}, /* 0x828c */
            {8'h00}, /* 0x828b */
            {8'h00}, /* 0x828a */
            {8'h00}, /* 0x8289 */
            {8'h00}, /* 0x8288 */
            {8'h00}, /* 0x8287 */
            {8'h00}, /* 0x8286 */
            {8'h00}, /* 0x8285 */
            {8'h00}, /* 0x8284 */
            {8'h00}, /* 0x8283 */
            {8'h00}, /* 0x8282 */
            {8'h00}, /* 0x8281 */
            {8'h00}, /* 0x8280 */
            {8'h00}, /* 0x827f */
            {8'h00}, /* 0x827e */
            {8'h00}, /* 0x827d */
            {8'h00}, /* 0x827c */
            {8'h00}, /* 0x827b */
            {8'h00}, /* 0x827a */
            {8'h00}, /* 0x8279 */
            {8'h00}, /* 0x8278 */
            {8'h00}, /* 0x8277 */
            {8'h00}, /* 0x8276 */
            {8'h00}, /* 0x8275 */
            {8'h00}, /* 0x8274 */
            {8'h00}, /* 0x8273 */
            {8'h00}, /* 0x8272 */
            {8'h00}, /* 0x8271 */
            {8'h00}, /* 0x8270 */
            {8'h00}, /* 0x826f */
            {8'h00}, /* 0x826e */
            {8'h00}, /* 0x826d */
            {8'h00}, /* 0x826c */
            {8'h00}, /* 0x826b */
            {8'h00}, /* 0x826a */
            {8'h00}, /* 0x8269 */
            {8'h00}, /* 0x8268 */
            {8'h00}, /* 0x8267 */
            {8'h00}, /* 0x8266 */
            {8'h00}, /* 0x8265 */
            {8'h00}, /* 0x8264 */
            {8'h00}, /* 0x8263 */
            {8'h00}, /* 0x8262 */
            {8'h00}, /* 0x8261 */
            {8'h00}, /* 0x8260 */
            {8'h00}, /* 0x825f */
            {8'h00}, /* 0x825e */
            {8'h00}, /* 0x825d */
            {8'h00}, /* 0x825c */
            {8'h00}, /* 0x825b */
            {8'h00}, /* 0x825a */
            {8'h00}, /* 0x8259 */
            {8'h00}, /* 0x8258 */
            {8'h00}, /* 0x8257 */
            {8'h00}, /* 0x8256 */
            {8'h00}, /* 0x8255 */
            {8'h00}, /* 0x8254 */
            {8'h00}, /* 0x8253 */
            {8'h00}, /* 0x8252 */
            {8'h00}, /* 0x8251 */
            {8'h00}, /* 0x8250 */
            {8'h00}, /* 0x824f */
            {8'h00}, /* 0x824e */
            {8'h00}, /* 0x824d */
            {8'h00}, /* 0x824c */
            {8'h00}, /* 0x824b */
            {8'h00}, /* 0x824a */
            {8'h00}, /* 0x8249 */
            {8'h00}, /* 0x8248 */
            {8'h00}, /* 0x8247 */
            {8'h00}, /* 0x8246 */
            {8'h00}, /* 0x8245 */
            {8'h00}, /* 0x8244 */
            {8'h00}, /* 0x8243 */
            {8'h00}, /* 0x8242 */
            {8'h00}, /* 0x8241 */
            {8'h00}, /* 0x8240 */
            {8'h00}, /* 0x823f */
            {8'h00}, /* 0x823e */
            {8'h00}, /* 0x823d */
            {8'h00}, /* 0x823c */
            {8'h00}, /* 0x823b */
            {8'h00}, /* 0x823a */
            {8'h00}, /* 0x8239 */
            {8'h00}, /* 0x8238 */
            {8'h00}, /* 0x8237 */
            {8'h00}, /* 0x8236 */
            {8'h00}, /* 0x8235 */
            {8'h00}, /* 0x8234 */
            {8'h00}, /* 0x8233 */
            {8'h00}, /* 0x8232 */
            {8'h00}, /* 0x8231 */
            {8'h00}, /* 0x8230 */
            {8'h00}, /* 0x822f */
            {8'h00}, /* 0x822e */
            {8'h00}, /* 0x822d */
            {8'h00}, /* 0x822c */
            {8'h00}, /* 0x822b */
            {8'h00}, /* 0x822a */
            {8'h00}, /* 0x8229 */
            {8'h00}, /* 0x8228 */
            {8'h00}, /* 0x8227 */
            {8'h00}, /* 0x8226 */
            {8'h00}, /* 0x8225 */
            {8'h00}, /* 0x8224 */
            {8'h00}, /* 0x8223 */
            {8'h00}, /* 0x8222 */
            {8'h00}, /* 0x8221 */
            {8'h00}, /* 0x8220 */
            {8'h00}, /* 0x821f */
            {8'h00}, /* 0x821e */
            {8'h00}, /* 0x821d */
            {8'h00}, /* 0x821c */
            {8'h00}, /* 0x821b */
            {8'h00}, /* 0x821a */
            {8'h00}, /* 0x8219 */
            {8'h00}, /* 0x8218 */
            {8'h00}, /* 0x8217 */
            {8'h00}, /* 0x8216 */
            {8'h00}, /* 0x8215 */
            {8'h00}, /* 0x8214 */
            {8'h00}, /* 0x8213 */
            {8'h00}, /* 0x8212 */
            {8'h00}, /* 0x8211 */
            {8'h00}, /* 0x8210 */
            {8'h00}, /* 0x820f */
            {8'h00}, /* 0x820e */
            {8'h00}, /* 0x820d */
            {8'h00}, /* 0x820c */
            {8'h00}, /* 0x820b */
            {8'h00}, /* 0x820a */
            {8'h00}, /* 0x8209 */
            {8'h00}, /* 0x8208 */
            {8'h00}, /* 0x8207 */
            {8'h00}, /* 0x8206 */
            {8'h00}, /* 0x8205 */
            {8'h00}, /* 0x8204 */
            {8'h00}, /* 0x8203 */
            {8'h00}, /* 0x8202 */
            {8'h00}, /* 0x8201 */
            {8'h00}, /* 0x8200 */
            {8'h00}, /* 0x81ff */
            {8'h00}, /* 0x81fe */
            {8'h00}, /* 0x81fd */
            {8'h00}, /* 0x81fc */
            {8'h00}, /* 0x81fb */
            {8'h00}, /* 0x81fa */
            {8'h00}, /* 0x81f9 */
            {8'h00}, /* 0x81f8 */
            {8'h00}, /* 0x81f7 */
            {8'h00}, /* 0x81f6 */
            {8'h00}, /* 0x81f5 */
            {8'h00}, /* 0x81f4 */
            {8'h00}, /* 0x81f3 */
            {8'h00}, /* 0x81f2 */
            {8'h00}, /* 0x81f1 */
            {8'h00}, /* 0x81f0 */
            {8'h00}, /* 0x81ef */
            {8'h00}, /* 0x81ee */
            {8'h00}, /* 0x81ed */
            {8'h00}, /* 0x81ec */
            {8'h00}, /* 0x81eb */
            {8'h00}, /* 0x81ea */
            {8'h00}, /* 0x81e9 */
            {8'h00}, /* 0x81e8 */
            {8'h00}, /* 0x81e7 */
            {8'h00}, /* 0x81e6 */
            {8'h00}, /* 0x81e5 */
            {8'h00}, /* 0x81e4 */
            {8'h00}, /* 0x81e3 */
            {8'h00}, /* 0x81e2 */
            {8'h00}, /* 0x81e1 */
            {8'h00}, /* 0x81e0 */
            {8'h00}, /* 0x81df */
            {8'h00}, /* 0x81de */
            {8'h00}, /* 0x81dd */
            {8'h00}, /* 0x81dc */
            {8'h00}, /* 0x81db */
            {8'h00}, /* 0x81da */
            {8'h00}, /* 0x81d9 */
            {8'h00}, /* 0x81d8 */
            {8'h00}, /* 0x81d7 */
            {8'h00}, /* 0x81d6 */
            {8'h00}, /* 0x81d5 */
            {8'h00}, /* 0x81d4 */
            {8'h00}, /* 0x81d3 */
            {8'h00}, /* 0x81d2 */
            {8'h00}, /* 0x81d1 */
            {8'h00}, /* 0x81d0 */
            {8'h00}, /* 0x81cf */
            {8'h00}, /* 0x81ce */
            {8'h00}, /* 0x81cd */
            {8'h00}, /* 0x81cc */
            {8'h00}, /* 0x81cb */
            {8'h00}, /* 0x81ca */
            {8'h00}, /* 0x81c9 */
            {8'h00}, /* 0x81c8 */
            {8'h00}, /* 0x81c7 */
            {8'h00}, /* 0x81c6 */
            {8'h00}, /* 0x81c5 */
            {8'h00}, /* 0x81c4 */
            {8'h00}, /* 0x81c3 */
            {8'h00}, /* 0x81c2 */
            {8'h00}, /* 0x81c1 */
            {8'h00}, /* 0x81c0 */
            {8'h00}, /* 0x81bf */
            {8'h00}, /* 0x81be */
            {8'h00}, /* 0x81bd */
            {8'h00}, /* 0x81bc */
            {8'h00}, /* 0x81bb */
            {8'h00}, /* 0x81ba */
            {8'h00}, /* 0x81b9 */
            {8'h00}, /* 0x81b8 */
            {8'h00}, /* 0x81b7 */
            {8'h00}, /* 0x81b6 */
            {8'h00}, /* 0x81b5 */
            {8'h00}, /* 0x81b4 */
            {8'h00}, /* 0x81b3 */
            {8'h00}, /* 0x81b2 */
            {8'h00}, /* 0x81b1 */
            {8'h00}, /* 0x81b0 */
            {8'h00}, /* 0x81af */
            {8'h00}, /* 0x81ae */
            {8'h00}, /* 0x81ad */
            {8'h00}, /* 0x81ac */
            {8'h00}, /* 0x81ab */
            {8'h00}, /* 0x81aa */
            {8'h00}, /* 0x81a9 */
            {8'h00}, /* 0x81a8 */
            {8'h00}, /* 0x81a7 */
            {8'h00}, /* 0x81a6 */
            {8'h00}, /* 0x81a5 */
            {8'h00}, /* 0x81a4 */
            {8'h00}, /* 0x81a3 */
            {8'h00}, /* 0x81a2 */
            {8'h00}, /* 0x81a1 */
            {8'h00}, /* 0x81a0 */
            {8'h00}, /* 0x819f */
            {8'h00}, /* 0x819e */
            {8'h00}, /* 0x819d */
            {8'h00}, /* 0x819c */
            {8'h00}, /* 0x819b */
            {8'h00}, /* 0x819a */
            {8'h00}, /* 0x8199 */
            {8'h00}, /* 0x8198 */
            {8'h00}, /* 0x8197 */
            {8'h00}, /* 0x8196 */
            {8'h00}, /* 0x8195 */
            {8'h00}, /* 0x8194 */
            {8'h00}, /* 0x8193 */
            {8'h00}, /* 0x8192 */
            {8'h00}, /* 0x8191 */
            {8'h00}, /* 0x8190 */
            {8'h00}, /* 0x818f */
            {8'h00}, /* 0x818e */
            {8'h00}, /* 0x818d */
            {8'h00}, /* 0x818c */
            {8'h00}, /* 0x818b */
            {8'h00}, /* 0x818a */
            {8'h00}, /* 0x8189 */
            {8'h00}, /* 0x8188 */
            {8'h00}, /* 0x8187 */
            {8'h00}, /* 0x8186 */
            {8'h00}, /* 0x8185 */
            {8'h00}, /* 0x8184 */
            {8'h00}, /* 0x8183 */
            {8'h00}, /* 0x8182 */
            {8'h00}, /* 0x8181 */
            {8'h00}, /* 0x8180 */
            {8'h00}, /* 0x817f */
            {8'h00}, /* 0x817e */
            {8'h00}, /* 0x817d */
            {8'h00}, /* 0x817c */
            {8'h00}, /* 0x817b */
            {8'h00}, /* 0x817a */
            {8'h00}, /* 0x8179 */
            {8'h00}, /* 0x8178 */
            {8'h00}, /* 0x8177 */
            {8'h00}, /* 0x8176 */
            {8'h00}, /* 0x8175 */
            {8'h00}, /* 0x8174 */
            {8'h00}, /* 0x8173 */
            {8'h00}, /* 0x8172 */
            {8'h00}, /* 0x8171 */
            {8'h00}, /* 0x8170 */
            {8'h00}, /* 0x816f */
            {8'h00}, /* 0x816e */
            {8'h00}, /* 0x816d */
            {8'h00}, /* 0x816c */
            {8'h00}, /* 0x816b */
            {8'h00}, /* 0x816a */
            {8'h00}, /* 0x8169 */
            {8'h00}, /* 0x8168 */
            {8'h00}, /* 0x8167 */
            {8'h00}, /* 0x8166 */
            {8'h00}, /* 0x8165 */
            {8'h00}, /* 0x8164 */
            {8'h00}, /* 0x8163 */
            {8'h00}, /* 0x8162 */
            {8'h00}, /* 0x8161 */
            {8'h00}, /* 0x8160 */
            {8'h00}, /* 0x815f */
            {8'h00}, /* 0x815e */
            {8'h00}, /* 0x815d */
            {8'h00}, /* 0x815c */
            {8'h00}, /* 0x815b */
            {8'h00}, /* 0x815a */
            {8'h00}, /* 0x8159 */
            {8'h00}, /* 0x8158 */
            {8'h00}, /* 0x8157 */
            {8'h00}, /* 0x8156 */
            {8'h00}, /* 0x8155 */
            {8'h00}, /* 0x8154 */
            {8'h00}, /* 0x8153 */
            {8'h00}, /* 0x8152 */
            {8'h00}, /* 0x8151 */
            {8'h00}, /* 0x8150 */
            {8'h00}, /* 0x814f */
            {8'h00}, /* 0x814e */
            {8'h00}, /* 0x814d */
            {8'h00}, /* 0x814c */
            {8'h00}, /* 0x814b */
            {8'h00}, /* 0x814a */
            {8'h00}, /* 0x8149 */
            {8'h00}, /* 0x8148 */
            {8'h00}, /* 0x8147 */
            {8'h00}, /* 0x8146 */
            {8'h00}, /* 0x8145 */
            {8'h00}, /* 0x8144 */
            {8'h00}, /* 0x8143 */
            {8'h00}, /* 0x8142 */
            {8'h00}, /* 0x8141 */
            {8'h00}, /* 0x8140 */
            {8'h00}, /* 0x813f */
            {8'h00}, /* 0x813e */
            {8'h00}, /* 0x813d */
            {8'h00}, /* 0x813c */
            {8'h00}, /* 0x813b */
            {8'h00}, /* 0x813a */
            {8'h00}, /* 0x8139 */
            {8'h00}, /* 0x8138 */
            {8'h00}, /* 0x8137 */
            {8'h00}, /* 0x8136 */
            {8'h00}, /* 0x8135 */
            {8'h00}, /* 0x8134 */
            {8'h00}, /* 0x8133 */
            {8'h00}, /* 0x8132 */
            {8'h00}, /* 0x8131 */
            {8'h00}, /* 0x8130 */
            {8'h00}, /* 0x812f */
            {8'h00}, /* 0x812e */
            {8'h00}, /* 0x812d */
            {8'h00}, /* 0x812c */
            {8'h00}, /* 0x812b */
            {8'h00}, /* 0x812a */
            {8'h00}, /* 0x8129 */
            {8'h00}, /* 0x8128 */
            {8'h00}, /* 0x8127 */
            {8'h00}, /* 0x8126 */
            {8'h00}, /* 0x8125 */
            {8'h00}, /* 0x8124 */
            {8'h00}, /* 0x8123 */
            {8'h00}, /* 0x8122 */
            {8'h00}, /* 0x8121 */
            {8'h00}, /* 0x8120 */
            {8'h00}, /* 0x811f */
            {8'h00}, /* 0x811e */
            {8'h00}, /* 0x811d */
            {8'h00}, /* 0x811c */
            {8'h00}, /* 0x811b */
            {8'h00}, /* 0x811a */
            {8'h00}, /* 0x8119 */
            {8'h00}, /* 0x8118 */
            {8'h00}, /* 0x8117 */
            {8'h00}, /* 0x8116 */
            {8'h00}, /* 0x8115 */
            {8'h00}, /* 0x8114 */
            {8'h00}, /* 0x8113 */
            {8'h00}, /* 0x8112 */
            {8'h00}, /* 0x8111 */
            {8'h00}, /* 0x8110 */
            {8'h00}, /* 0x810f */
            {8'h00}, /* 0x810e */
            {8'h00}, /* 0x810d */
            {8'h00}, /* 0x810c */
            {8'h00}, /* 0x810b */
            {8'h00}, /* 0x810a */
            {8'h00}, /* 0x8109 */
            {8'h00}, /* 0x8108 */
            {8'h00}, /* 0x8107 */
            {8'h00}, /* 0x8106 */
            {8'h00}, /* 0x8105 */
            {8'h00}, /* 0x8104 */
            {8'h00}, /* 0x8103 */
            {8'h00}, /* 0x8102 */
            {8'h00}, /* 0x8101 */
            {8'h00}, /* 0x8100 */
            {8'h00}, /* 0x80ff */
            {8'h00}, /* 0x80fe */
            {8'h00}, /* 0x80fd */
            {8'h00}, /* 0x80fc */
            {8'h00}, /* 0x80fb */
            {8'h00}, /* 0x80fa */
            {8'h00}, /* 0x80f9 */
            {8'h00}, /* 0x80f8 */
            {8'h00}, /* 0x80f7 */
            {8'h00}, /* 0x80f6 */
            {8'h00}, /* 0x80f5 */
            {8'h00}, /* 0x80f4 */
            {8'h00}, /* 0x80f3 */
            {8'h00}, /* 0x80f2 */
            {8'h00}, /* 0x80f1 */
            {8'h00}, /* 0x80f0 */
            {8'h00}, /* 0x80ef */
            {8'h00}, /* 0x80ee */
            {8'h00}, /* 0x80ed */
            {8'h00}, /* 0x80ec */
            {8'h00}, /* 0x80eb */
            {8'h00}, /* 0x80ea */
            {8'h00}, /* 0x80e9 */
            {8'h00}, /* 0x80e8 */
            {8'h00}, /* 0x80e7 */
            {8'h00}, /* 0x80e6 */
            {8'h00}, /* 0x80e5 */
            {8'h00}, /* 0x80e4 */
            {8'h00}, /* 0x80e3 */
            {8'h00}, /* 0x80e2 */
            {8'h00}, /* 0x80e1 */
            {8'h00}, /* 0x80e0 */
            {8'h00}, /* 0x80df */
            {8'h00}, /* 0x80de */
            {8'h00}, /* 0x80dd */
            {8'h00}, /* 0x80dc */
            {8'h00}, /* 0x80db */
            {8'h00}, /* 0x80da */
            {8'h00}, /* 0x80d9 */
            {8'h00}, /* 0x80d8 */
            {8'h00}, /* 0x80d7 */
            {8'h00}, /* 0x80d6 */
            {8'h00}, /* 0x80d5 */
            {8'h00}, /* 0x80d4 */
            {8'h00}, /* 0x80d3 */
            {8'h00}, /* 0x80d2 */
            {8'h00}, /* 0x80d1 */
            {8'h00}, /* 0x80d0 */
            {8'h00}, /* 0x80cf */
            {8'h00}, /* 0x80ce */
            {8'h00}, /* 0x80cd */
            {8'h00}, /* 0x80cc */
            {8'h00}, /* 0x80cb */
            {8'h00}, /* 0x80ca */
            {8'h00}, /* 0x80c9 */
            {8'h00}, /* 0x80c8 */
            {8'h00}, /* 0x80c7 */
            {8'h00}, /* 0x80c6 */
            {8'h00}, /* 0x80c5 */
            {8'h00}, /* 0x80c4 */
            {8'h00}, /* 0x80c3 */
            {8'h00}, /* 0x80c2 */
            {8'h00}, /* 0x80c1 */
            {8'h00}, /* 0x80c0 */
            {8'h00}, /* 0x80bf */
            {8'h00}, /* 0x80be */
            {8'h00}, /* 0x80bd */
            {8'h00}, /* 0x80bc */
            {8'h00}, /* 0x80bb */
            {8'h00}, /* 0x80ba */
            {8'h00}, /* 0x80b9 */
            {8'h00}, /* 0x80b8 */
            {8'h00}, /* 0x80b7 */
            {8'h00}, /* 0x80b6 */
            {8'h00}, /* 0x80b5 */
            {8'h00}, /* 0x80b4 */
            {8'h00}, /* 0x80b3 */
            {8'h00}, /* 0x80b2 */
            {8'h00}, /* 0x80b1 */
            {8'h00}, /* 0x80b0 */
            {8'h00}, /* 0x80af */
            {8'h00}, /* 0x80ae */
            {8'h00}, /* 0x80ad */
            {8'h00}, /* 0x80ac */
            {8'h00}, /* 0x80ab */
            {8'h00}, /* 0x80aa */
            {8'h00}, /* 0x80a9 */
            {8'h00}, /* 0x80a8 */
            {8'h00}, /* 0x80a7 */
            {8'h00}, /* 0x80a6 */
            {8'h00}, /* 0x80a5 */
            {8'h00}, /* 0x80a4 */
            {8'h00}, /* 0x80a3 */
            {8'h00}, /* 0x80a2 */
            {8'h00}, /* 0x80a1 */
            {8'h00}, /* 0x80a0 */
            {8'h00}, /* 0x809f */
            {8'h00}, /* 0x809e */
            {8'h00}, /* 0x809d */
            {8'h00}, /* 0x809c */
            {8'h00}, /* 0x809b */
            {8'h00}, /* 0x809a */
            {8'h00}, /* 0x8099 */
            {8'h00}, /* 0x8098 */
            {8'h00}, /* 0x8097 */
            {8'h00}, /* 0x8096 */
            {8'h00}, /* 0x8095 */
            {8'h00}, /* 0x8094 */
            {8'h00}, /* 0x8093 */
            {8'h00}, /* 0x8092 */
            {8'h00}, /* 0x8091 */
            {8'h00}, /* 0x8090 */
            {8'h00}, /* 0x808f */
            {8'h00}, /* 0x808e */
            {8'h00}, /* 0x808d */
            {8'h00}, /* 0x808c */
            {8'h00}, /* 0x808b */
            {8'h00}, /* 0x808a */
            {8'h00}, /* 0x8089 */
            {8'h00}, /* 0x8088 */
            {8'h00}, /* 0x8087 */
            {8'h00}, /* 0x8086 */
            {8'h00}, /* 0x8085 */
            {8'h00}, /* 0x8084 */
            {8'h00}, /* 0x8083 */
            {8'h00}, /* 0x8082 */
            {8'h00}, /* 0x8081 */
            {8'h00}, /* 0x8080 */
            {8'h00}, /* 0x807f */
            {8'h00}, /* 0x807e */
            {8'h00}, /* 0x807d */
            {8'h00}, /* 0x807c */
            {8'h00}, /* 0x807b */
            {8'h00}, /* 0x807a */
            {8'h00}, /* 0x8079 */
            {8'h00}, /* 0x8078 */
            {8'h00}, /* 0x8077 */
            {8'h00}, /* 0x8076 */
            {8'h00}, /* 0x8075 */
            {8'h00}, /* 0x8074 */
            {8'h00}, /* 0x8073 */
            {8'h00}, /* 0x8072 */
            {8'h00}, /* 0x8071 */
            {8'h00}, /* 0x8070 */
            {8'h00}, /* 0x806f */
            {8'h00}, /* 0x806e */
            {8'h00}, /* 0x806d */
            {8'h00}, /* 0x806c */
            {8'h00}, /* 0x806b */
            {8'h00}, /* 0x806a */
            {8'h00}, /* 0x8069 */
            {8'h00}, /* 0x8068 */
            {8'h00}, /* 0x8067 */
            {8'h00}, /* 0x8066 */
            {8'h00}, /* 0x8065 */
            {8'h00}, /* 0x8064 */
            {8'h00}, /* 0x8063 */
            {8'h00}, /* 0x8062 */
            {8'h00}, /* 0x8061 */
            {8'h00}, /* 0x8060 */
            {8'h00}, /* 0x805f */
            {8'h00}, /* 0x805e */
            {8'h00}, /* 0x805d */
            {8'h00}, /* 0x805c */
            {8'h00}, /* 0x805b */
            {8'h00}, /* 0x805a */
            {8'h00}, /* 0x8059 */
            {8'h00}, /* 0x8058 */
            {8'h00}, /* 0x8057 */
            {8'h00}, /* 0x8056 */
            {8'h00}, /* 0x8055 */
            {8'h00}, /* 0x8054 */
            {8'h00}, /* 0x8053 */
            {8'h00}, /* 0x8052 */
            {8'h00}, /* 0x8051 */
            {8'h00}, /* 0x8050 */
            {8'h00}, /* 0x804f */
            {8'h00}, /* 0x804e */
            {8'h00}, /* 0x804d */
            {8'h00}, /* 0x804c */
            {8'h00}, /* 0x804b */
            {8'h00}, /* 0x804a */
            {8'h00}, /* 0x8049 */
            {8'h00}, /* 0x8048 */
            {8'h00}, /* 0x8047 */
            {8'h00}, /* 0x8046 */
            {8'h00}, /* 0x8045 */
            {8'h00}, /* 0x8044 */
            {8'h00}, /* 0x8043 */
            {8'h00}, /* 0x8042 */
            {8'h00}, /* 0x8041 */
            {8'h00}, /* 0x8040 */
            {8'h00}, /* 0x803f */
            {8'h00}, /* 0x803e */
            {8'h00}, /* 0x803d */
            {8'h00}, /* 0x803c */
            {8'h00}, /* 0x803b */
            {8'h00}, /* 0x803a */
            {8'h00}, /* 0x8039 */
            {8'h00}, /* 0x8038 */
            {8'h00}, /* 0x8037 */
            {8'h00}, /* 0x8036 */
            {8'h00}, /* 0x8035 */
            {8'h00}, /* 0x8034 */
            {8'h00}, /* 0x8033 */
            {8'h00}, /* 0x8032 */
            {8'h00}, /* 0x8031 */
            {8'h00}, /* 0x8030 */
            {8'h00}, /* 0x802f */
            {8'h00}, /* 0x802e */
            {8'h00}, /* 0x802d */
            {8'h00}, /* 0x802c */
            {8'h00}, /* 0x802b */
            {8'h00}, /* 0x802a */
            {8'h00}, /* 0x8029 */
            {8'h00}, /* 0x8028 */
            {8'h00}, /* 0x8027 */
            {8'h00}, /* 0x8026 */
            {8'h00}, /* 0x8025 */
            {8'h00}, /* 0x8024 */
            {8'h00}, /* 0x8023 */
            {8'h00}, /* 0x8022 */
            {8'h00}, /* 0x8021 */
            {8'h00}, /* 0x8020 */
            {8'h00}, /* 0x801f */
            {8'h00}, /* 0x801e */
            {8'h00}, /* 0x801d */
            {8'h00}, /* 0x801c */
            {8'h00}, /* 0x801b */
            {8'h00}, /* 0x801a */
            {8'h00}, /* 0x8019 */
            {8'h00}, /* 0x8018 */
            {8'h00}, /* 0x8017 */
            {8'h00}, /* 0x8016 */
            {8'h00}, /* 0x8015 */
            {8'h00}, /* 0x8014 */
            {8'h00}, /* 0x8013 */
            {8'h00}, /* 0x8012 */
            {8'h00}, /* 0x8011 */
            {8'h00}, /* 0x8010 */
            {8'h00}, /* 0x800f */
            {8'h00}, /* 0x800e */
            {8'h00}, /* 0x800d */
            {8'h00}, /* 0x800c */
            {8'h00}, /* 0x800b */
            {8'h00}, /* 0x800a */
            {8'h00}, /* 0x8009 */
            {8'h00}, /* 0x8008 */
            {8'h00}, /* 0x8007 */
            {8'h00}, /* 0x8006 */
            {8'h00}, /* 0x8005 */
            {8'h00}, /* 0x8004 */
            {8'h00}, /* 0x8003 */
            {8'h00}, /* 0x8002 */
            {8'h00}, /* 0x8001 */
            {8'h00}, /* 0x8000 */
            {8'h00}, /* 0x7fff */
            {8'h00}, /* 0x7ffe */
            {8'h00}, /* 0x7ffd */
            {8'h00}, /* 0x7ffc */
            {8'h00}, /* 0x7ffb */
            {8'h00}, /* 0x7ffa */
            {8'h00}, /* 0x7ff9 */
            {8'h00}, /* 0x7ff8 */
            {8'h00}, /* 0x7ff7 */
            {8'h00}, /* 0x7ff6 */
            {8'h00}, /* 0x7ff5 */
            {8'h00}, /* 0x7ff4 */
            {8'h00}, /* 0x7ff3 */
            {8'h00}, /* 0x7ff2 */
            {8'h00}, /* 0x7ff1 */
            {8'h00}, /* 0x7ff0 */
            {8'h00}, /* 0x7fef */
            {8'h00}, /* 0x7fee */
            {8'h00}, /* 0x7fed */
            {8'h00}, /* 0x7fec */
            {8'h00}, /* 0x7feb */
            {8'h00}, /* 0x7fea */
            {8'h00}, /* 0x7fe9 */
            {8'h00}, /* 0x7fe8 */
            {8'h00}, /* 0x7fe7 */
            {8'h00}, /* 0x7fe6 */
            {8'h00}, /* 0x7fe5 */
            {8'h00}, /* 0x7fe4 */
            {8'h00}, /* 0x7fe3 */
            {8'h00}, /* 0x7fe2 */
            {8'h00}, /* 0x7fe1 */
            {8'h00}, /* 0x7fe0 */
            {8'h00}, /* 0x7fdf */
            {8'h00}, /* 0x7fde */
            {8'h00}, /* 0x7fdd */
            {8'h00}, /* 0x7fdc */
            {8'h00}, /* 0x7fdb */
            {8'h00}, /* 0x7fda */
            {8'h00}, /* 0x7fd9 */
            {8'h00}, /* 0x7fd8 */
            {8'h00}, /* 0x7fd7 */
            {8'h00}, /* 0x7fd6 */
            {8'h00}, /* 0x7fd5 */
            {8'h00}, /* 0x7fd4 */
            {8'h00}, /* 0x7fd3 */
            {8'h00}, /* 0x7fd2 */
            {8'h00}, /* 0x7fd1 */
            {8'h00}, /* 0x7fd0 */
            {8'h00}, /* 0x7fcf */
            {8'h00}, /* 0x7fce */
            {8'h00}, /* 0x7fcd */
            {8'h00}, /* 0x7fcc */
            {8'h00}, /* 0x7fcb */
            {8'h00}, /* 0x7fca */
            {8'h00}, /* 0x7fc9 */
            {8'h00}, /* 0x7fc8 */
            {8'h00}, /* 0x7fc7 */
            {8'h00}, /* 0x7fc6 */
            {8'h00}, /* 0x7fc5 */
            {8'h00}, /* 0x7fc4 */
            {8'h00}, /* 0x7fc3 */
            {8'h00}, /* 0x7fc2 */
            {8'h00}, /* 0x7fc1 */
            {8'h00}, /* 0x7fc0 */
            {8'h00}, /* 0x7fbf */
            {8'h00}, /* 0x7fbe */
            {8'h00}, /* 0x7fbd */
            {8'h00}, /* 0x7fbc */
            {8'h00}, /* 0x7fbb */
            {8'h00}, /* 0x7fba */
            {8'h00}, /* 0x7fb9 */
            {8'h00}, /* 0x7fb8 */
            {8'h00}, /* 0x7fb7 */
            {8'h00}, /* 0x7fb6 */
            {8'h00}, /* 0x7fb5 */
            {8'h00}, /* 0x7fb4 */
            {8'h00}, /* 0x7fb3 */
            {8'h00}, /* 0x7fb2 */
            {8'h00}, /* 0x7fb1 */
            {8'h00}, /* 0x7fb0 */
            {8'h00}, /* 0x7faf */
            {8'h00}, /* 0x7fae */
            {8'h00}, /* 0x7fad */
            {8'h00}, /* 0x7fac */
            {8'h00}, /* 0x7fab */
            {8'h00}, /* 0x7faa */
            {8'h00}, /* 0x7fa9 */
            {8'h00}, /* 0x7fa8 */
            {8'h00}, /* 0x7fa7 */
            {8'h00}, /* 0x7fa6 */
            {8'h00}, /* 0x7fa5 */
            {8'h00}, /* 0x7fa4 */
            {8'h00}, /* 0x7fa3 */
            {8'h00}, /* 0x7fa2 */
            {8'h00}, /* 0x7fa1 */
            {8'h00}, /* 0x7fa0 */
            {8'h00}, /* 0x7f9f */
            {8'h00}, /* 0x7f9e */
            {8'h00}, /* 0x7f9d */
            {8'h00}, /* 0x7f9c */
            {8'h00}, /* 0x7f9b */
            {8'h00}, /* 0x7f9a */
            {8'h00}, /* 0x7f99 */
            {8'h00}, /* 0x7f98 */
            {8'h00}, /* 0x7f97 */
            {8'h00}, /* 0x7f96 */
            {8'h00}, /* 0x7f95 */
            {8'h00}, /* 0x7f94 */
            {8'h00}, /* 0x7f93 */
            {8'h00}, /* 0x7f92 */
            {8'h00}, /* 0x7f91 */
            {8'h00}, /* 0x7f90 */
            {8'h00}, /* 0x7f8f */
            {8'h00}, /* 0x7f8e */
            {8'h00}, /* 0x7f8d */
            {8'h00}, /* 0x7f8c */
            {8'h00}, /* 0x7f8b */
            {8'h00}, /* 0x7f8a */
            {8'h00}, /* 0x7f89 */
            {8'h00}, /* 0x7f88 */
            {8'h00}, /* 0x7f87 */
            {8'h00}, /* 0x7f86 */
            {8'h00}, /* 0x7f85 */
            {8'h00}, /* 0x7f84 */
            {8'h00}, /* 0x7f83 */
            {8'h00}, /* 0x7f82 */
            {8'h00}, /* 0x7f81 */
            {8'h00}, /* 0x7f80 */
            {8'h00}, /* 0x7f7f */
            {8'h00}, /* 0x7f7e */
            {8'h00}, /* 0x7f7d */
            {8'h00}, /* 0x7f7c */
            {8'h00}, /* 0x7f7b */
            {8'h00}, /* 0x7f7a */
            {8'h00}, /* 0x7f79 */
            {8'h00}, /* 0x7f78 */
            {8'h00}, /* 0x7f77 */
            {8'h00}, /* 0x7f76 */
            {8'h00}, /* 0x7f75 */
            {8'h00}, /* 0x7f74 */
            {8'h00}, /* 0x7f73 */
            {8'h00}, /* 0x7f72 */
            {8'h00}, /* 0x7f71 */
            {8'h00}, /* 0x7f70 */
            {8'h00}, /* 0x7f6f */
            {8'h00}, /* 0x7f6e */
            {8'h00}, /* 0x7f6d */
            {8'h00}, /* 0x7f6c */
            {8'h00}, /* 0x7f6b */
            {8'h00}, /* 0x7f6a */
            {8'h00}, /* 0x7f69 */
            {8'h00}, /* 0x7f68 */
            {8'h00}, /* 0x7f67 */
            {8'h00}, /* 0x7f66 */
            {8'h00}, /* 0x7f65 */
            {8'h00}, /* 0x7f64 */
            {8'h00}, /* 0x7f63 */
            {8'h00}, /* 0x7f62 */
            {8'h00}, /* 0x7f61 */
            {8'h00}, /* 0x7f60 */
            {8'h00}, /* 0x7f5f */
            {8'h00}, /* 0x7f5e */
            {8'h00}, /* 0x7f5d */
            {8'h00}, /* 0x7f5c */
            {8'h00}, /* 0x7f5b */
            {8'h00}, /* 0x7f5a */
            {8'h00}, /* 0x7f59 */
            {8'h00}, /* 0x7f58 */
            {8'h00}, /* 0x7f57 */
            {8'h00}, /* 0x7f56 */
            {8'h00}, /* 0x7f55 */
            {8'h00}, /* 0x7f54 */
            {8'h00}, /* 0x7f53 */
            {8'h00}, /* 0x7f52 */
            {8'h00}, /* 0x7f51 */
            {8'h00}, /* 0x7f50 */
            {8'h00}, /* 0x7f4f */
            {8'h00}, /* 0x7f4e */
            {8'h00}, /* 0x7f4d */
            {8'h00}, /* 0x7f4c */
            {8'h00}, /* 0x7f4b */
            {8'h00}, /* 0x7f4a */
            {8'h00}, /* 0x7f49 */
            {8'h00}, /* 0x7f48 */
            {8'h00}, /* 0x7f47 */
            {8'h00}, /* 0x7f46 */
            {8'h00}, /* 0x7f45 */
            {8'h00}, /* 0x7f44 */
            {8'h00}, /* 0x7f43 */
            {8'h00}, /* 0x7f42 */
            {8'h00}, /* 0x7f41 */
            {8'h00}, /* 0x7f40 */
            {8'h00}, /* 0x7f3f */
            {8'h00}, /* 0x7f3e */
            {8'h00}, /* 0x7f3d */
            {8'h00}, /* 0x7f3c */
            {8'h00}, /* 0x7f3b */
            {8'h00}, /* 0x7f3a */
            {8'h00}, /* 0x7f39 */
            {8'h00}, /* 0x7f38 */
            {8'h00}, /* 0x7f37 */
            {8'h00}, /* 0x7f36 */
            {8'h00}, /* 0x7f35 */
            {8'h00}, /* 0x7f34 */
            {8'h00}, /* 0x7f33 */
            {8'h00}, /* 0x7f32 */
            {8'h00}, /* 0x7f31 */
            {8'h00}, /* 0x7f30 */
            {8'h00}, /* 0x7f2f */
            {8'h00}, /* 0x7f2e */
            {8'h00}, /* 0x7f2d */
            {8'h00}, /* 0x7f2c */
            {8'h00}, /* 0x7f2b */
            {8'h00}, /* 0x7f2a */
            {8'h00}, /* 0x7f29 */
            {8'h00}, /* 0x7f28 */
            {8'h00}, /* 0x7f27 */
            {8'h00}, /* 0x7f26 */
            {8'h00}, /* 0x7f25 */
            {8'h00}, /* 0x7f24 */
            {8'h00}, /* 0x7f23 */
            {8'h00}, /* 0x7f22 */
            {8'h00}, /* 0x7f21 */
            {8'h00}, /* 0x7f20 */
            {8'h00}, /* 0x7f1f */
            {8'h00}, /* 0x7f1e */
            {8'h00}, /* 0x7f1d */
            {8'h00}, /* 0x7f1c */
            {8'h00}, /* 0x7f1b */
            {8'h00}, /* 0x7f1a */
            {8'h00}, /* 0x7f19 */
            {8'h00}, /* 0x7f18 */
            {8'h00}, /* 0x7f17 */
            {8'h00}, /* 0x7f16 */
            {8'h00}, /* 0x7f15 */
            {8'h00}, /* 0x7f14 */
            {8'h00}, /* 0x7f13 */
            {8'h00}, /* 0x7f12 */
            {8'h00}, /* 0x7f11 */
            {8'h00}, /* 0x7f10 */
            {8'h00}, /* 0x7f0f */
            {8'h00}, /* 0x7f0e */
            {8'h00}, /* 0x7f0d */
            {8'h00}, /* 0x7f0c */
            {8'h00}, /* 0x7f0b */
            {8'h00}, /* 0x7f0a */
            {8'h00}, /* 0x7f09 */
            {8'h00}, /* 0x7f08 */
            {8'h00}, /* 0x7f07 */
            {8'h00}, /* 0x7f06 */
            {8'h00}, /* 0x7f05 */
            {8'h00}, /* 0x7f04 */
            {8'h00}, /* 0x7f03 */
            {8'h00}, /* 0x7f02 */
            {8'h00}, /* 0x7f01 */
            {8'h00}, /* 0x7f00 */
            {8'h00}, /* 0x7eff */
            {8'h00}, /* 0x7efe */
            {8'h00}, /* 0x7efd */
            {8'h00}, /* 0x7efc */
            {8'h00}, /* 0x7efb */
            {8'h00}, /* 0x7efa */
            {8'h00}, /* 0x7ef9 */
            {8'h00}, /* 0x7ef8 */
            {8'h00}, /* 0x7ef7 */
            {8'h00}, /* 0x7ef6 */
            {8'h00}, /* 0x7ef5 */
            {8'h00}, /* 0x7ef4 */
            {8'h00}, /* 0x7ef3 */
            {8'h00}, /* 0x7ef2 */
            {8'h00}, /* 0x7ef1 */
            {8'h00}, /* 0x7ef0 */
            {8'h00}, /* 0x7eef */
            {8'h00}, /* 0x7eee */
            {8'h00}, /* 0x7eed */
            {8'h00}, /* 0x7eec */
            {8'h00}, /* 0x7eeb */
            {8'h00}, /* 0x7eea */
            {8'h00}, /* 0x7ee9 */
            {8'h00}, /* 0x7ee8 */
            {8'h00}, /* 0x7ee7 */
            {8'h00}, /* 0x7ee6 */
            {8'h00}, /* 0x7ee5 */
            {8'h00}, /* 0x7ee4 */
            {8'h00}, /* 0x7ee3 */
            {8'h00}, /* 0x7ee2 */
            {8'h00}, /* 0x7ee1 */
            {8'h00}, /* 0x7ee0 */
            {8'h00}, /* 0x7edf */
            {8'h00}, /* 0x7ede */
            {8'h00}, /* 0x7edd */
            {8'h00}, /* 0x7edc */
            {8'h00}, /* 0x7edb */
            {8'h00}, /* 0x7eda */
            {8'h00}, /* 0x7ed9 */
            {8'h00}, /* 0x7ed8 */
            {8'h00}, /* 0x7ed7 */
            {8'h00}, /* 0x7ed6 */
            {8'h00}, /* 0x7ed5 */
            {8'h00}, /* 0x7ed4 */
            {8'h00}, /* 0x7ed3 */
            {8'h00}, /* 0x7ed2 */
            {8'h00}, /* 0x7ed1 */
            {8'h00}, /* 0x7ed0 */
            {8'h00}, /* 0x7ecf */
            {8'h00}, /* 0x7ece */
            {8'h00}, /* 0x7ecd */
            {8'h00}, /* 0x7ecc */
            {8'h00}, /* 0x7ecb */
            {8'h00}, /* 0x7eca */
            {8'h00}, /* 0x7ec9 */
            {8'h00}, /* 0x7ec8 */
            {8'h00}, /* 0x7ec7 */
            {8'h00}, /* 0x7ec6 */
            {8'h00}, /* 0x7ec5 */
            {8'h00}, /* 0x7ec4 */
            {8'h00}, /* 0x7ec3 */
            {8'h00}, /* 0x7ec2 */
            {8'h00}, /* 0x7ec1 */
            {8'h00}, /* 0x7ec0 */
            {8'h00}, /* 0x7ebf */
            {8'h00}, /* 0x7ebe */
            {8'h00}, /* 0x7ebd */
            {8'h00}, /* 0x7ebc */
            {8'h00}, /* 0x7ebb */
            {8'h00}, /* 0x7eba */
            {8'h00}, /* 0x7eb9 */
            {8'h00}, /* 0x7eb8 */
            {8'h00}, /* 0x7eb7 */
            {8'h00}, /* 0x7eb6 */
            {8'h00}, /* 0x7eb5 */
            {8'h00}, /* 0x7eb4 */
            {8'h00}, /* 0x7eb3 */
            {8'h00}, /* 0x7eb2 */
            {8'h00}, /* 0x7eb1 */
            {8'h00}, /* 0x7eb0 */
            {8'h00}, /* 0x7eaf */
            {8'h00}, /* 0x7eae */
            {8'h00}, /* 0x7ead */
            {8'h00}, /* 0x7eac */
            {8'h00}, /* 0x7eab */
            {8'h00}, /* 0x7eaa */
            {8'h00}, /* 0x7ea9 */
            {8'h00}, /* 0x7ea8 */
            {8'h00}, /* 0x7ea7 */
            {8'h00}, /* 0x7ea6 */
            {8'h00}, /* 0x7ea5 */
            {8'h00}, /* 0x7ea4 */
            {8'h00}, /* 0x7ea3 */
            {8'h00}, /* 0x7ea2 */
            {8'h00}, /* 0x7ea1 */
            {8'h00}, /* 0x7ea0 */
            {8'h00}, /* 0x7e9f */
            {8'h00}, /* 0x7e9e */
            {8'h00}, /* 0x7e9d */
            {8'h00}, /* 0x7e9c */
            {8'h00}, /* 0x7e9b */
            {8'h00}, /* 0x7e9a */
            {8'h00}, /* 0x7e99 */
            {8'h00}, /* 0x7e98 */
            {8'h00}, /* 0x7e97 */
            {8'h00}, /* 0x7e96 */
            {8'h00}, /* 0x7e95 */
            {8'h00}, /* 0x7e94 */
            {8'h00}, /* 0x7e93 */
            {8'h00}, /* 0x7e92 */
            {8'h00}, /* 0x7e91 */
            {8'h00}, /* 0x7e90 */
            {8'h00}, /* 0x7e8f */
            {8'h00}, /* 0x7e8e */
            {8'h00}, /* 0x7e8d */
            {8'h00}, /* 0x7e8c */
            {8'h00}, /* 0x7e8b */
            {8'h00}, /* 0x7e8a */
            {8'h00}, /* 0x7e89 */
            {8'h00}, /* 0x7e88 */
            {8'h00}, /* 0x7e87 */
            {8'h00}, /* 0x7e86 */
            {8'h00}, /* 0x7e85 */
            {8'h00}, /* 0x7e84 */
            {8'h00}, /* 0x7e83 */
            {8'h00}, /* 0x7e82 */
            {8'h00}, /* 0x7e81 */
            {8'h00}, /* 0x7e80 */
            {8'h00}, /* 0x7e7f */
            {8'h00}, /* 0x7e7e */
            {8'h00}, /* 0x7e7d */
            {8'h00}, /* 0x7e7c */
            {8'h00}, /* 0x7e7b */
            {8'h00}, /* 0x7e7a */
            {8'h00}, /* 0x7e79 */
            {8'h00}, /* 0x7e78 */
            {8'h00}, /* 0x7e77 */
            {8'h00}, /* 0x7e76 */
            {8'h00}, /* 0x7e75 */
            {8'h00}, /* 0x7e74 */
            {8'h00}, /* 0x7e73 */
            {8'h00}, /* 0x7e72 */
            {8'h00}, /* 0x7e71 */
            {8'h00}, /* 0x7e70 */
            {8'h00}, /* 0x7e6f */
            {8'h00}, /* 0x7e6e */
            {8'h00}, /* 0x7e6d */
            {8'h00}, /* 0x7e6c */
            {8'h00}, /* 0x7e6b */
            {8'h00}, /* 0x7e6a */
            {8'h00}, /* 0x7e69 */
            {8'h00}, /* 0x7e68 */
            {8'h00}, /* 0x7e67 */
            {8'h00}, /* 0x7e66 */
            {8'h00}, /* 0x7e65 */
            {8'h00}, /* 0x7e64 */
            {8'h00}, /* 0x7e63 */
            {8'h00}, /* 0x7e62 */
            {8'h00}, /* 0x7e61 */
            {8'h00}, /* 0x7e60 */
            {8'h00}, /* 0x7e5f */
            {8'h00}, /* 0x7e5e */
            {8'h00}, /* 0x7e5d */
            {8'h00}, /* 0x7e5c */
            {8'h00}, /* 0x7e5b */
            {8'h00}, /* 0x7e5a */
            {8'h00}, /* 0x7e59 */
            {8'h00}, /* 0x7e58 */
            {8'h00}, /* 0x7e57 */
            {8'h00}, /* 0x7e56 */
            {8'h00}, /* 0x7e55 */
            {8'h00}, /* 0x7e54 */
            {8'h00}, /* 0x7e53 */
            {8'h00}, /* 0x7e52 */
            {8'h00}, /* 0x7e51 */
            {8'h00}, /* 0x7e50 */
            {8'h00}, /* 0x7e4f */
            {8'h00}, /* 0x7e4e */
            {8'h00}, /* 0x7e4d */
            {8'h00}, /* 0x7e4c */
            {8'h00}, /* 0x7e4b */
            {8'h00}, /* 0x7e4a */
            {8'h00}, /* 0x7e49 */
            {8'h00}, /* 0x7e48 */
            {8'h00}, /* 0x7e47 */
            {8'h00}, /* 0x7e46 */
            {8'h00}, /* 0x7e45 */
            {8'h00}, /* 0x7e44 */
            {8'h00}, /* 0x7e43 */
            {8'h00}, /* 0x7e42 */
            {8'h00}, /* 0x7e41 */
            {8'h00}, /* 0x7e40 */
            {8'h00}, /* 0x7e3f */
            {8'h00}, /* 0x7e3e */
            {8'h00}, /* 0x7e3d */
            {8'h00}, /* 0x7e3c */
            {8'h00}, /* 0x7e3b */
            {8'h00}, /* 0x7e3a */
            {8'h00}, /* 0x7e39 */
            {8'h00}, /* 0x7e38 */
            {8'h00}, /* 0x7e37 */
            {8'h00}, /* 0x7e36 */
            {8'h00}, /* 0x7e35 */
            {8'h00}, /* 0x7e34 */
            {8'h00}, /* 0x7e33 */
            {8'h00}, /* 0x7e32 */
            {8'h00}, /* 0x7e31 */
            {8'h00}, /* 0x7e30 */
            {8'h00}, /* 0x7e2f */
            {8'h00}, /* 0x7e2e */
            {8'h00}, /* 0x7e2d */
            {8'h00}, /* 0x7e2c */
            {8'h00}, /* 0x7e2b */
            {8'h00}, /* 0x7e2a */
            {8'h00}, /* 0x7e29 */
            {8'h00}, /* 0x7e28 */
            {8'h00}, /* 0x7e27 */
            {8'h00}, /* 0x7e26 */
            {8'h00}, /* 0x7e25 */
            {8'h00}, /* 0x7e24 */
            {8'h00}, /* 0x7e23 */
            {8'h00}, /* 0x7e22 */
            {8'h00}, /* 0x7e21 */
            {8'h00}, /* 0x7e20 */
            {8'h00}, /* 0x7e1f */
            {8'h00}, /* 0x7e1e */
            {8'h00}, /* 0x7e1d */
            {8'h00}, /* 0x7e1c */
            {8'h00}, /* 0x7e1b */
            {8'h00}, /* 0x7e1a */
            {8'h00}, /* 0x7e19 */
            {8'h00}, /* 0x7e18 */
            {8'h00}, /* 0x7e17 */
            {8'h00}, /* 0x7e16 */
            {8'h00}, /* 0x7e15 */
            {8'h00}, /* 0x7e14 */
            {8'h00}, /* 0x7e13 */
            {8'h00}, /* 0x7e12 */
            {8'h00}, /* 0x7e11 */
            {8'h00}, /* 0x7e10 */
            {8'h00}, /* 0x7e0f */
            {8'h00}, /* 0x7e0e */
            {8'h00}, /* 0x7e0d */
            {8'h00}, /* 0x7e0c */
            {8'h00}, /* 0x7e0b */
            {8'h00}, /* 0x7e0a */
            {8'h00}, /* 0x7e09 */
            {8'h00}, /* 0x7e08 */
            {8'h00}, /* 0x7e07 */
            {8'h00}, /* 0x7e06 */
            {8'h00}, /* 0x7e05 */
            {8'h00}, /* 0x7e04 */
            {8'h00}, /* 0x7e03 */
            {8'h00}, /* 0x7e02 */
            {8'h00}, /* 0x7e01 */
            {8'h00}, /* 0x7e00 */
            {8'h00}, /* 0x7dff */
            {8'h00}, /* 0x7dfe */
            {8'h00}, /* 0x7dfd */
            {8'h00}, /* 0x7dfc */
            {8'h00}, /* 0x7dfb */
            {8'h00}, /* 0x7dfa */
            {8'h00}, /* 0x7df9 */
            {8'h00}, /* 0x7df8 */
            {8'h00}, /* 0x7df7 */
            {8'h00}, /* 0x7df6 */
            {8'h00}, /* 0x7df5 */
            {8'h00}, /* 0x7df4 */
            {8'h00}, /* 0x7df3 */
            {8'h00}, /* 0x7df2 */
            {8'h00}, /* 0x7df1 */
            {8'h00}, /* 0x7df0 */
            {8'h00}, /* 0x7def */
            {8'h00}, /* 0x7dee */
            {8'h00}, /* 0x7ded */
            {8'h00}, /* 0x7dec */
            {8'h00}, /* 0x7deb */
            {8'h00}, /* 0x7dea */
            {8'h00}, /* 0x7de9 */
            {8'h00}, /* 0x7de8 */
            {8'h00}, /* 0x7de7 */
            {8'h00}, /* 0x7de6 */
            {8'h00}, /* 0x7de5 */
            {8'h00}, /* 0x7de4 */
            {8'h00}, /* 0x7de3 */
            {8'h00}, /* 0x7de2 */
            {8'h00}, /* 0x7de1 */
            {8'h00}, /* 0x7de0 */
            {8'h00}, /* 0x7ddf */
            {8'h00}, /* 0x7dde */
            {8'h00}, /* 0x7ddd */
            {8'h00}, /* 0x7ddc */
            {8'h00}, /* 0x7ddb */
            {8'h00}, /* 0x7dda */
            {8'h00}, /* 0x7dd9 */
            {8'h00}, /* 0x7dd8 */
            {8'h00}, /* 0x7dd7 */
            {8'h00}, /* 0x7dd6 */
            {8'h00}, /* 0x7dd5 */
            {8'h00}, /* 0x7dd4 */
            {8'h00}, /* 0x7dd3 */
            {8'h00}, /* 0x7dd2 */
            {8'h00}, /* 0x7dd1 */
            {8'h00}, /* 0x7dd0 */
            {8'h00}, /* 0x7dcf */
            {8'h00}, /* 0x7dce */
            {8'h00}, /* 0x7dcd */
            {8'h00}, /* 0x7dcc */
            {8'h00}, /* 0x7dcb */
            {8'h00}, /* 0x7dca */
            {8'h00}, /* 0x7dc9 */
            {8'h00}, /* 0x7dc8 */
            {8'h00}, /* 0x7dc7 */
            {8'h00}, /* 0x7dc6 */
            {8'h00}, /* 0x7dc5 */
            {8'h00}, /* 0x7dc4 */
            {8'h00}, /* 0x7dc3 */
            {8'h00}, /* 0x7dc2 */
            {8'h00}, /* 0x7dc1 */
            {8'h00}, /* 0x7dc0 */
            {8'h00}, /* 0x7dbf */
            {8'h00}, /* 0x7dbe */
            {8'h00}, /* 0x7dbd */
            {8'h00}, /* 0x7dbc */
            {8'h00}, /* 0x7dbb */
            {8'h00}, /* 0x7dba */
            {8'h00}, /* 0x7db9 */
            {8'h00}, /* 0x7db8 */
            {8'h00}, /* 0x7db7 */
            {8'h00}, /* 0x7db6 */
            {8'h00}, /* 0x7db5 */
            {8'h00}, /* 0x7db4 */
            {8'h00}, /* 0x7db3 */
            {8'h00}, /* 0x7db2 */
            {8'h00}, /* 0x7db1 */
            {8'h00}, /* 0x7db0 */
            {8'h00}, /* 0x7daf */
            {8'h00}, /* 0x7dae */
            {8'h00}, /* 0x7dad */
            {8'h00}, /* 0x7dac */
            {8'h00}, /* 0x7dab */
            {8'h00}, /* 0x7daa */
            {8'h00}, /* 0x7da9 */
            {8'h00}, /* 0x7da8 */
            {8'h00}, /* 0x7da7 */
            {8'h00}, /* 0x7da6 */
            {8'h00}, /* 0x7da5 */
            {8'h00}, /* 0x7da4 */
            {8'h00}, /* 0x7da3 */
            {8'h00}, /* 0x7da2 */
            {8'h00}, /* 0x7da1 */
            {8'h00}, /* 0x7da0 */
            {8'h00}, /* 0x7d9f */
            {8'h00}, /* 0x7d9e */
            {8'h00}, /* 0x7d9d */
            {8'h00}, /* 0x7d9c */
            {8'h00}, /* 0x7d9b */
            {8'h00}, /* 0x7d9a */
            {8'h00}, /* 0x7d99 */
            {8'h00}, /* 0x7d98 */
            {8'h00}, /* 0x7d97 */
            {8'h00}, /* 0x7d96 */
            {8'h00}, /* 0x7d95 */
            {8'h00}, /* 0x7d94 */
            {8'h00}, /* 0x7d93 */
            {8'h00}, /* 0x7d92 */
            {8'h00}, /* 0x7d91 */
            {8'h00}, /* 0x7d90 */
            {8'h00}, /* 0x7d8f */
            {8'h00}, /* 0x7d8e */
            {8'h00}, /* 0x7d8d */
            {8'h00}, /* 0x7d8c */
            {8'h00}, /* 0x7d8b */
            {8'h00}, /* 0x7d8a */
            {8'h00}, /* 0x7d89 */
            {8'h00}, /* 0x7d88 */
            {8'h00}, /* 0x7d87 */
            {8'h00}, /* 0x7d86 */
            {8'h00}, /* 0x7d85 */
            {8'h00}, /* 0x7d84 */
            {8'h00}, /* 0x7d83 */
            {8'h00}, /* 0x7d82 */
            {8'h00}, /* 0x7d81 */
            {8'h00}, /* 0x7d80 */
            {8'h00}, /* 0x7d7f */
            {8'h00}, /* 0x7d7e */
            {8'h00}, /* 0x7d7d */
            {8'h00}, /* 0x7d7c */
            {8'h00}, /* 0x7d7b */
            {8'h00}, /* 0x7d7a */
            {8'h00}, /* 0x7d79 */
            {8'h00}, /* 0x7d78 */
            {8'h00}, /* 0x7d77 */
            {8'h00}, /* 0x7d76 */
            {8'h00}, /* 0x7d75 */
            {8'h00}, /* 0x7d74 */
            {8'h00}, /* 0x7d73 */
            {8'h00}, /* 0x7d72 */
            {8'h00}, /* 0x7d71 */
            {8'h00}, /* 0x7d70 */
            {8'h00}, /* 0x7d6f */
            {8'h00}, /* 0x7d6e */
            {8'h00}, /* 0x7d6d */
            {8'h00}, /* 0x7d6c */
            {8'h00}, /* 0x7d6b */
            {8'h00}, /* 0x7d6a */
            {8'h00}, /* 0x7d69 */
            {8'h00}, /* 0x7d68 */
            {8'h00}, /* 0x7d67 */
            {8'h00}, /* 0x7d66 */
            {8'h00}, /* 0x7d65 */
            {8'h00}, /* 0x7d64 */
            {8'h00}, /* 0x7d63 */
            {8'h00}, /* 0x7d62 */
            {8'h00}, /* 0x7d61 */
            {8'h00}, /* 0x7d60 */
            {8'h00}, /* 0x7d5f */
            {8'h00}, /* 0x7d5e */
            {8'h00}, /* 0x7d5d */
            {8'h00}, /* 0x7d5c */
            {8'h00}, /* 0x7d5b */
            {8'h00}, /* 0x7d5a */
            {8'h00}, /* 0x7d59 */
            {8'h00}, /* 0x7d58 */
            {8'h00}, /* 0x7d57 */
            {8'h00}, /* 0x7d56 */
            {8'h00}, /* 0x7d55 */
            {8'h00}, /* 0x7d54 */
            {8'h00}, /* 0x7d53 */
            {8'h00}, /* 0x7d52 */
            {8'h00}, /* 0x7d51 */
            {8'h00}, /* 0x7d50 */
            {8'h00}, /* 0x7d4f */
            {8'h00}, /* 0x7d4e */
            {8'h00}, /* 0x7d4d */
            {8'h00}, /* 0x7d4c */
            {8'h00}, /* 0x7d4b */
            {8'h00}, /* 0x7d4a */
            {8'h00}, /* 0x7d49 */
            {8'h00}, /* 0x7d48 */
            {8'h00}, /* 0x7d47 */
            {8'h00}, /* 0x7d46 */
            {8'h00}, /* 0x7d45 */
            {8'h00}, /* 0x7d44 */
            {8'h00}, /* 0x7d43 */
            {8'h00}, /* 0x7d42 */
            {8'h00}, /* 0x7d41 */
            {8'h00}, /* 0x7d40 */
            {8'h00}, /* 0x7d3f */
            {8'h00}, /* 0x7d3e */
            {8'h00}, /* 0x7d3d */
            {8'h00}, /* 0x7d3c */
            {8'h00}, /* 0x7d3b */
            {8'h00}, /* 0x7d3a */
            {8'h00}, /* 0x7d39 */
            {8'h00}, /* 0x7d38 */
            {8'h00}, /* 0x7d37 */
            {8'h00}, /* 0x7d36 */
            {8'h00}, /* 0x7d35 */
            {8'h00}, /* 0x7d34 */
            {8'h00}, /* 0x7d33 */
            {8'h00}, /* 0x7d32 */
            {8'h00}, /* 0x7d31 */
            {8'h00}, /* 0x7d30 */
            {8'h00}, /* 0x7d2f */
            {8'h00}, /* 0x7d2e */
            {8'h00}, /* 0x7d2d */
            {8'h00}, /* 0x7d2c */
            {8'h00}, /* 0x7d2b */
            {8'h00}, /* 0x7d2a */
            {8'h00}, /* 0x7d29 */
            {8'h00}, /* 0x7d28 */
            {8'h00}, /* 0x7d27 */
            {8'h00}, /* 0x7d26 */
            {8'h00}, /* 0x7d25 */
            {8'h00}, /* 0x7d24 */
            {8'h00}, /* 0x7d23 */
            {8'h00}, /* 0x7d22 */
            {8'h00}, /* 0x7d21 */
            {8'h00}, /* 0x7d20 */
            {8'h00}, /* 0x7d1f */
            {8'h00}, /* 0x7d1e */
            {8'h00}, /* 0x7d1d */
            {8'h00}, /* 0x7d1c */
            {8'h00}, /* 0x7d1b */
            {8'h00}, /* 0x7d1a */
            {8'h00}, /* 0x7d19 */
            {8'h00}, /* 0x7d18 */
            {8'h00}, /* 0x7d17 */
            {8'h00}, /* 0x7d16 */
            {8'h00}, /* 0x7d15 */
            {8'h00}, /* 0x7d14 */
            {8'h00}, /* 0x7d13 */
            {8'h00}, /* 0x7d12 */
            {8'h00}, /* 0x7d11 */
            {8'h00}, /* 0x7d10 */
            {8'h00}, /* 0x7d0f */
            {8'h00}, /* 0x7d0e */
            {8'h00}, /* 0x7d0d */
            {8'h00}, /* 0x7d0c */
            {8'h00}, /* 0x7d0b */
            {8'h00}, /* 0x7d0a */
            {8'h00}, /* 0x7d09 */
            {8'h00}, /* 0x7d08 */
            {8'h00}, /* 0x7d07 */
            {8'h00}, /* 0x7d06 */
            {8'h00}, /* 0x7d05 */
            {8'h00}, /* 0x7d04 */
            {8'h00}, /* 0x7d03 */
            {8'h00}, /* 0x7d02 */
            {8'h00}, /* 0x7d01 */
            {8'h00}, /* 0x7d00 */
            {8'h00}, /* 0x7cff */
            {8'h00}, /* 0x7cfe */
            {8'h00}, /* 0x7cfd */
            {8'h00}, /* 0x7cfc */
            {8'h00}, /* 0x7cfb */
            {8'h00}, /* 0x7cfa */
            {8'h00}, /* 0x7cf9 */
            {8'h00}, /* 0x7cf8 */
            {8'h00}, /* 0x7cf7 */
            {8'h00}, /* 0x7cf6 */
            {8'h00}, /* 0x7cf5 */
            {8'h00}, /* 0x7cf4 */
            {8'h00}, /* 0x7cf3 */
            {8'h00}, /* 0x7cf2 */
            {8'h00}, /* 0x7cf1 */
            {8'h00}, /* 0x7cf0 */
            {8'h00}, /* 0x7cef */
            {8'h00}, /* 0x7cee */
            {8'h00}, /* 0x7ced */
            {8'h00}, /* 0x7cec */
            {8'h00}, /* 0x7ceb */
            {8'h00}, /* 0x7cea */
            {8'h00}, /* 0x7ce9 */
            {8'h00}, /* 0x7ce8 */
            {8'h00}, /* 0x7ce7 */
            {8'h00}, /* 0x7ce6 */
            {8'h00}, /* 0x7ce5 */
            {8'h00}, /* 0x7ce4 */
            {8'h00}, /* 0x7ce3 */
            {8'h00}, /* 0x7ce2 */
            {8'h00}, /* 0x7ce1 */
            {8'h00}, /* 0x7ce0 */
            {8'h00}, /* 0x7cdf */
            {8'h00}, /* 0x7cde */
            {8'h00}, /* 0x7cdd */
            {8'h00}, /* 0x7cdc */
            {8'h00}, /* 0x7cdb */
            {8'h00}, /* 0x7cda */
            {8'h00}, /* 0x7cd9 */
            {8'h00}, /* 0x7cd8 */
            {8'h00}, /* 0x7cd7 */
            {8'h00}, /* 0x7cd6 */
            {8'h00}, /* 0x7cd5 */
            {8'h00}, /* 0x7cd4 */
            {8'h00}, /* 0x7cd3 */
            {8'h00}, /* 0x7cd2 */
            {8'h00}, /* 0x7cd1 */
            {8'h00}, /* 0x7cd0 */
            {8'h00}, /* 0x7ccf */
            {8'h00}, /* 0x7cce */
            {8'h00}, /* 0x7ccd */
            {8'h00}, /* 0x7ccc */
            {8'h00}, /* 0x7ccb */
            {8'h00}, /* 0x7cca */
            {8'h00}, /* 0x7cc9 */
            {8'h00}, /* 0x7cc8 */
            {8'h00}, /* 0x7cc7 */
            {8'h00}, /* 0x7cc6 */
            {8'h00}, /* 0x7cc5 */
            {8'h00}, /* 0x7cc4 */
            {8'h00}, /* 0x7cc3 */
            {8'h00}, /* 0x7cc2 */
            {8'h00}, /* 0x7cc1 */
            {8'h00}, /* 0x7cc0 */
            {8'h00}, /* 0x7cbf */
            {8'h00}, /* 0x7cbe */
            {8'h00}, /* 0x7cbd */
            {8'h00}, /* 0x7cbc */
            {8'h00}, /* 0x7cbb */
            {8'h00}, /* 0x7cba */
            {8'h00}, /* 0x7cb9 */
            {8'h00}, /* 0x7cb8 */
            {8'h00}, /* 0x7cb7 */
            {8'h00}, /* 0x7cb6 */
            {8'h00}, /* 0x7cb5 */
            {8'h00}, /* 0x7cb4 */
            {8'h00}, /* 0x7cb3 */
            {8'h00}, /* 0x7cb2 */
            {8'h00}, /* 0x7cb1 */
            {8'h00}, /* 0x7cb0 */
            {8'h00}, /* 0x7caf */
            {8'h00}, /* 0x7cae */
            {8'h00}, /* 0x7cad */
            {8'h00}, /* 0x7cac */
            {8'h00}, /* 0x7cab */
            {8'h00}, /* 0x7caa */
            {8'h00}, /* 0x7ca9 */
            {8'h00}, /* 0x7ca8 */
            {8'h00}, /* 0x7ca7 */
            {8'h00}, /* 0x7ca6 */
            {8'h00}, /* 0x7ca5 */
            {8'h00}, /* 0x7ca4 */
            {8'h00}, /* 0x7ca3 */
            {8'h00}, /* 0x7ca2 */
            {8'h00}, /* 0x7ca1 */
            {8'h00}, /* 0x7ca0 */
            {8'h00}, /* 0x7c9f */
            {8'h00}, /* 0x7c9e */
            {8'h00}, /* 0x7c9d */
            {8'h00}, /* 0x7c9c */
            {8'h00}, /* 0x7c9b */
            {8'h00}, /* 0x7c9a */
            {8'h00}, /* 0x7c99 */
            {8'h00}, /* 0x7c98 */
            {8'h00}, /* 0x7c97 */
            {8'h00}, /* 0x7c96 */
            {8'h00}, /* 0x7c95 */
            {8'h00}, /* 0x7c94 */
            {8'h00}, /* 0x7c93 */
            {8'h00}, /* 0x7c92 */
            {8'h00}, /* 0x7c91 */
            {8'h00}, /* 0x7c90 */
            {8'h00}, /* 0x7c8f */
            {8'h00}, /* 0x7c8e */
            {8'h00}, /* 0x7c8d */
            {8'h00}, /* 0x7c8c */
            {8'h00}, /* 0x7c8b */
            {8'h00}, /* 0x7c8a */
            {8'h00}, /* 0x7c89 */
            {8'h00}, /* 0x7c88 */
            {8'h00}, /* 0x7c87 */
            {8'h00}, /* 0x7c86 */
            {8'h00}, /* 0x7c85 */
            {8'h00}, /* 0x7c84 */
            {8'h00}, /* 0x7c83 */
            {8'h00}, /* 0x7c82 */
            {8'h00}, /* 0x7c81 */
            {8'h00}, /* 0x7c80 */
            {8'h00}, /* 0x7c7f */
            {8'h00}, /* 0x7c7e */
            {8'h00}, /* 0x7c7d */
            {8'h00}, /* 0x7c7c */
            {8'h00}, /* 0x7c7b */
            {8'h00}, /* 0x7c7a */
            {8'h00}, /* 0x7c79 */
            {8'h00}, /* 0x7c78 */
            {8'h00}, /* 0x7c77 */
            {8'h00}, /* 0x7c76 */
            {8'h00}, /* 0x7c75 */
            {8'h00}, /* 0x7c74 */
            {8'h00}, /* 0x7c73 */
            {8'h00}, /* 0x7c72 */
            {8'h00}, /* 0x7c71 */
            {8'h00}, /* 0x7c70 */
            {8'h00}, /* 0x7c6f */
            {8'h00}, /* 0x7c6e */
            {8'h00}, /* 0x7c6d */
            {8'h00}, /* 0x7c6c */
            {8'h00}, /* 0x7c6b */
            {8'h00}, /* 0x7c6a */
            {8'h00}, /* 0x7c69 */
            {8'h00}, /* 0x7c68 */
            {8'h00}, /* 0x7c67 */
            {8'h00}, /* 0x7c66 */
            {8'h00}, /* 0x7c65 */
            {8'h00}, /* 0x7c64 */
            {8'h00}, /* 0x7c63 */
            {8'h00}, /* 0x7c62 */
            {8'h00}, /* 0x7c61 */
            {8'h00}, /* 0x7c60 */
            {8'h00}, /* 0x7c5f */
            {8'h00}, /* 0x7c5e */
            {8'h00}, /* 0x7c5d */
            {8'h00}, /* 0x7c5c */
            {8'h00}, /* 0x7c5b */
            {8'h00}, /* 0x7c5a */
            {8'h00}, /* 0x7c59 */
            {8'h00}, /* 0x7c58 */
            {8'h00}, /* 0x7c57 */
            {8'h00}, /* 0x7c56 */
            {8'h00}, /* 0x7c55 */
            {8'h00}, /* 0x7c54 */
            {8'h00}, /* 0x7c53 */
            {8'h00}, /* 0x7c52 */
            {8'h00}, /* 0x7c51 */
            {8'h00}, /* 0x7c50 */
            {8'h00}, /* 0x7c4f */
            {8'h00}, /* 0x7c4e */
            {8'h00}, /* 0x7c4d */
            {8'h00}, /* 0x7c4c */
            {8'h00}, /* 0x7c4b */
            {8'h00}, /* 0x7c4a */
            {8'h00}, /* 0x7c49 */
            {8'h00}, /* 0x7c48 */
            {8'h00}, /* 0x7c47 */
            {8'h00}, /* 0x7c46 */
            {8'h00}, /* 0x7c45 */
            {8'h00}, /* 0x7c44 */
            {8'h00}, /* 0x7c43 */
            {8'h00}, /* 0x7c42 */
            {8'h00}, /* 0x7c41 */
            {8'h00}, /* 0x7c40 */
            {8'h00}, /* 0x7c3f */
            {8'h00}, /* 0x7c3e */
            {8'h00}, /* 0x7c3d */
            {8'h00}, /* 0x7c3c */
            {8'h00}, /* 0x7c3b */
            {8'h00}, /* 0x7c3a */
            {8'h00}, /* 0x7c39 */
            {8'h00}, /* 0x7c38 */
            {8'h00}, /* 0x7c37 */
            {8'h00}, /* 0x7c36 */
            {8'h00}, /* 0x7c35 */
            {8'h00}, /* 0x7c34 */
            {8'h00}, /* 0x7c33 */
            {8'h00}, /* 0x7c32 */
            {8'h00}, /* 0x7c31 */
            {8'h00}, /* 0x7c30 */
            {8'h00}, /* 0x7c2f */
            {8'h00}, /* 0x7c2e */
            {8'h00}, /* 0x7c2d */
            {8'h00}, /* 0x7c2c */
            {8'h00}, /* 0x7c2b */
            {8'h00}, /* 0x7c2a */
            {8'h00}, /* 0x7c29 */
            {8'h00}, /* 0x7c28 */
            {8'h00}, /* 0x7c27 */
            {8'h00}, /* 0x7c26 */
            {8'h00}, /* 0x7c25 */
            {8'h00}, /* 0x7c24 */
            {8'h00}, /* 0x7c23 */
            {8'h00}, /* 0x7c22 */
            {8'h00}, /* 0x7c21 */
            {8'h00}, /* 0x7c20 */
            {8'h00}, /* 0x7c1f */
            {8'h00}, /* 0x7c1e */
            {8'h00}, /* 0x7c1d */
            {8'h00}, /* 0x7c1c */
            {8'h00}, /* 0x7c1b */
            {8'h00}, /* 0x7c1a */
            {8'h00}, /* 0x7c19 */
            {8'h00}, /* 0x7c18 */
            {8'h00}, /* 0x7c17 */
            {8'h00}, /* 0x7c16 */
            {8'h00}, /* 0x7c15 */
            {8'h00}, /* 0x7c14 */
            {8'h00}, /* 0x7c13 */
            {8'h00}, /* 0x7c12 */
            {8'h00}, /* 0x7c11 */
            {8'h00}, /* 0x7c10 */
            {8'h00}, /* 0x7c0f */
            {8'h00}, /* 0x7c0e */
            {8'h00}, /* 0x7c0d */
            {8'h00}, /* 0x7c0c */
            {8'h00}, /* 0x7c0b */
            {8'h00}, /* 0x7c0a */
            {8'h00}, /* 0x7c09 */
            {8'h00}, /* 0x7c08 */
            {8'h00}, /* 0x7c07 */
            {8'h00}, /* 0x7c06 */
            {8'h00}, /* 0x7c05 */
            {8'h00}, /* 0x7c04 */
            {8'h00}, /* 0x7c03 */
            {8'h00}, /* 0x7c02 */
            {8'h00}, /* 0x7c01 */
            {8'h00}, /* 0x7c00 */
            {8'h00}, /* 0x7bff */
            {8'h00}, /* 0x7bfe */
            {8'h00}, /* 0x7bfd */
            {8'h00}, /* 0x7bfc */
            {8'h00}, /* 0x7bfb */
            {8'h00}, /* 0x7bfa */
            {8'h00}, /* 0x7bf9 */
            {8'h00}, /* 0x7bf8 */
            {8'h00}, /* 0x7bf7 */
            {8'h00}, /* 0x7bf6 */
            {8'h00}, /* 0x7bf5 */
            {8'h00}, /* 0x7bf4 */
            {8'h00}, /* 0x7bf3 */
            {8'h00}, /* 0x7bf2 */
            {8'h00}, /* 0x7bf1 */
            {8'h00}, /* 0x7bf0 */
            {8'h00}, /* 0x7bef */
            {8'h00}, /* 0x7bee */
            {8'h00}, /* 0x7bed */
            {8'h00}, /* 0x7bec */
            {8'h00}, /* 0x7beb */
            {8'h00}, /* 0x7bea */
            {8'h00}, /* 0x7be9 */
            {8'h00}, /* 0x7be8 */
            {8'h00}, /* 0x7be7 */
            {8'h00}, /* 0x7be6 */
            {8'h00}, /* 0x7be5 */
            {8'h00}, /* 0x7be4 */
            {8'h00}, /* 0x7be3 */
            {8'h00}, /* 0x7be2 */
            {8'h00}, /* 0x7be1 */
            {8'h00}, /* 0x7be0 */
            {8'h00}, /* 0x7bdf */
            {8'h00}, /* 0x7bde */
            {8'h00}, /* 0x7bdd */
            {8'h00}, /* 0x7bdc */
            {8'h00}, /* 0x7bdb */
            {8'h00}, /* 0x7bda */
            {8'h00}, /* 0x7bd9 */
            {8'h00}, /* 0x7bd8 */
            {8'h00}, /* 0x7bd7 */
            {8'h00}, /* 0x7bd6 */
            {8'h00}, /* 0x7bd5 */
            {8'h00}, /* 0x7bd4 */
            {8'h00}, /* 0x7bd3 */
            {8'h00}, /* 0x7bd2 */
            {8'h00}, /* 0x7bd1 */
            {8'h00}, /* 0x7bd0 */
            {8'h00}, /* 0x7bcf */
            {8'h00}, /* 0x7bce */
            {8'h00}, /* 0x7bcd */
            {8'h00}, /* 0x7bcc */
            {8'h00}, /* 0x7bcb */
            {8'h00}, /* 0x7bca */
            {8'h00}, /* 0x7bc9 */
            {8'h00}, /* 0x7bc8 */
            {8'h00}, /* 0x7bc7 */
            {8'h00}, /* 0x7bc6 */
            {8'h00}, /* 0x7bc5 */
            {8'h00}, /* 0x7bc4 */
            {8'h00}, /* 0x7bc3 */
            {8'h00}, /* 0x7bc2 */
            {8'h00}, /* 0x7bc1 */
            {8'h00}, /* 0x7bc0 */
            {8'h00}, /* 0x7bbf */
            {8'h00}, /* 0x7bbe */
            {8'h00}, /* 0x7bbd */
            {8'h00}, /* 0x7bbc */
            {8'h00}, /* 0x7bbb */
            {8'h00}, /* 0x7bba */
            {8'h00}, /* 0x7bb9 */
            {8'h00}, /* 0x7bb8 */
            {8'h00}, /* 0x7bb7 */
            {8'h00}, /* 0x7bb6 */
            {8'h00}, /* 0x7bb5 */
            {8'h00}, /* 0x7bb4 */
            {8'h00}, /* 0x7bb3 */
            {8'h00}, /* 0x7bb2 */
            {8'h00}, /* 0x7bb1 */
            {8'h00}, /* 0x7bb0 */
            {8'h00}, /* 0x7baf */
            {8'h00}, /* 0x7bae */
            {8'h00}, /* 0x7bad */
            {8'h00}, /* 0x7bac */
            {8'h00}, /* 0x7bab */
            {8'h00}, /* 0x7baa */
            {8'h00}, /* 0x7ba9 */
            {8'h00}, /* 0x7ba8 */
            {8'h00}, /* 0x7ba7 */
            {8'h00}, /* 0x7ba6 */
            {8'h00}, /* 0x7ba5 */
            {8'h00}, /* 0x7ba4 */
            {8'h00}, /* 0x7ba3 */
            {8'h00}, /* 0x7ba2 */
            {8'h00}, /* 0x7ba1 */
            {8'h00}, /* 0x7ba0 */
            {8'h00}, /* 0x7b9f */
            {8'h00}, /* 0x7b9e */
            {8'h00}, /* 0x7b9d */
            {8'h00}, /* 0x7b9c */
            {8'h00}, /* 0x7b9b */
            {8'h00}, /* 0x7b9a */
            {8'h00}, /* 0x7b99 */
            {8'h00}, /* 0x7b98 */
            {8'h00}, /* 0x7b97 */
            {8'h00}, /* 0x7b96 */
            {8'h00}, /* 0x7b95 */
            {8'h00}, /* 0x7b94 */
            {8'h00}, /* 0x7b93 */
            {8'h00}, /* 0x7b92 */
            {8'h00}, /* 0x7b91 */
            {8'h00}, /* 0x7b90 */
            {8'h00}, /* 0x7b8f */
            {8'h00}, /* 0x7b8e */
            {8'h00}, /* 0x7b8d */
            {8'h00}, /* 0x7b8c */
            {8'h00}, /* 0x7b8b */
            {8'h00}, /* 0x7b8a */
            {8'h00}, /* 0x7b89 */
            {8'h00}, /* 0x7b88 */
            {8'h00}, /* 0x7b87 */
            {8'h00}, /* 0x7b86 */
            {8'h00}, /* 0x7b85 */
            {8'h00}, /* 0x7b84 */
            {8'h00}, /* 0x7b83 */
            {8'h00}, /* 0x7b82 */
            {8'h00}, /* 0x7b81 */
            {8'h00}, /* 0x7b80 */
            {8'h00}, /* 0x7b7f */
            {8'h00}, /* 0x7b7e */
            {8'h00}, /* 0x7b7d */
            {8'h00}, /* 0x7b7c */
            {8'h00}, /* 0x7b7b */
            {8'h00}, /* 0x7b7a */
            {8'h00}, /* 0x7b79 */
            {8'h00}, /* 0x7b78 */
            {8'h00}, /* 0x7b77 */
            {8'h00}, /* 0x7b76 */
            {8'h00}, /* 0x7b75 */
            {8'h00}, /* 0x7b74 */
            {8'h00}, /* 0x7b73 */
            {8'h00}, /* 0x7b72 */
            {8'h00}, /* 0x7b71 */
            {8'h00}, /* 0x7b70 */
            {8'h00}, /* 0x7b6f */
            {8'h00}, /* 0x7b6e */
            {8'h00}, /* 0x7b6d */
            {8'h00}, /* 0x7b6c */
            {8'h00}, /* 0x7b6b */
            {8'h00}, /* 0x7b6a */
            {8'h00}, /* 0x7b69 */
            {8'h00}, /* 0x7b68 */
            {8'h00}, /* 0x7b67 */
            {8'h00}, /* 0x7b66 */
            {8'h00}, /* 0x7b65 */
            {8'h00}, /* 0x7b64 */
            {8'h00}, /* 0x7b63 */
            {8'h00}, /* 0x7b62 */
            {8'h00}, /* 0x7b61 */
            {8'h00}, /* 0x7b60 */
            {8'h00}, /* 0x7b5f */
            {8'h00}, /* 0x7b5e */
            {8'h00}, /* 0x7b5d */
            {8'h00}, /* 0x7b5c */
            {8'h00}, /* 0x7b5b */
            {8'h00}, /* 0x7b5a */
            {8'h00}, /* 0x7b59 */
            {8'h00}, /* 0x7b58 */
            {8'h00}, /* 0x7b57 */
            {8'h00}, /* 0x7b56 */
            {8'h00}, /* 0x7b55 */
            {8'h00}, /* 0x7b54 */
            {8'h00}, /* 0x7b53 */
            {8'h00}, /* 0x7b52 */
            {8'h00}, /* 0x7b51 */
            {8'h00}, /* 0x7b50 */
            {8'h00}, /* 0x7b4f */
            {8'h00}, /* 0x7b4e */
            {8'h00}, /* 0x7b4d */
            {8'h00}, /* 0x7b4c */
            {8'h00}, /* 0x7b4b */
            {8'h00}, /* 0x7b4a */
            {8'h00}, /* 0x7b49 */
            {8'h00}, /* 0x7b48 */
            {8'h00}, /* 0x7b47 */
            {8'h00}, /* 0x7b46 */
            {8'h00}, /* 0x7b45 */
            {8'h00}, /* 0x7b44 */
            {8'h00}, /* 0x7b43 */
            {8'h00}, /* 0x7b42 */
            {8'h00}, /* 0x7b41 */
            {8'h00}, /* 0x7b40 */
            {8'h00}, /* 0x7b3f */
            {8'h00}, /* 0x7b3e */
            {8'h00}, /* 0x7b3d */
            {8'h00}, /* 0x7b3c */
            {8'h00}, /* 0x7b3b */
            {8'h00}, /* 0x7b3a */
            {8'h00}, /* 0x7b39 */
            {8'h00}, /* 0x7b38 */
            {8'h00}, /* 0x7b37 */
            {8'h00}, /* 0x7b36 */
            {8'h00}, /* 0x7b35 */
            {8'h00}, /* 0x7b34 */
            {8'h00}, /* 0x7b33 */
            {8'h00}, /* 0x7b32 */
            {8'h00}, /* 0x7b31 */
            {8'h00}, /* 0x7b30 */
            {8'h00}, /* 0x7b2f */
            {8'h00}, /* 0x7b2e */
            {8'h00}, /* 0x7b2d */
            {8'h00}, /* 0x7b2c */
            {8'h00}, /* 0x7b2b */
            {8'h00}, /* 0x7b2a */
            {8'h00}, /* 0x7b29 */
            {8'h00}, /* 0x7b28 */
            {8'h00}, /* 0x7b27 */
            {8'h00}, /* 0x7b26 */
            {8'h00}, /* 0x7b25 */
            {8'h00}, /* 0x7b24 */
            {8'h00}, /* 0x7b23 */
            {8'h00}, /* 0x7b22 */
            {8'h00}, /* 0x7b21 */
            {8'h00}, /* 0x7b20 */
            {8'h00}, /* 0x7b1f */
            {8'h00}, /* 0x7b1e */
            {8'h00}, /* 0x7b1d */
            {8'h00}, /* 0x7b1c */
            {8'h00}, /* 0x7b1b */
            {8'h00}, /* 0x7b1a */
            {8'h00}, /* 0x7b19 */
            {8'h00}, /* 0x7b18 */
            {8'h00}, /* 0x7b17 */
            {8'h00}, /* 0x7b16 */
            {8'h00}, /* 0x7b15 */
            {8'h00}, /* 0x7b14 */
            {8'h00}, /* 0x7b13 */
            {8'h00}, /* 0x7b12 */
            {8'h00}, /* 0x7b11 */
            {8'h00}, /* 0x7b10 */
            {8'h00}, /* 0x7b0f */
            {8'h00}, /* 0x7b0e */
            {8'h00}, /* 0x7b0d */
            {8'h00}, /* 0x7b0c */
            {8'h00}, /* 0x7b0b */
            {8'h00}, /* 0x7b0a */
            {8'h00}, /* 0x7b09 */
            {8'h00}, /* 0x7b08 */
            {8'h00}, /* 0x7b07 */
            {8'h00}, /* 0x7b06 */
            {8'h00}, /* 0x7b05 */
            {8'h00}, /* 0x7b04 */
            {8'h00}, /* 0x7b03 */
            {8'h00}, /* 0x7b02 */
            {8'h00}, /* 0x7b01 */
            {8'h00}, /* 0x7b00 */
            {8'h00}, /* 0x7aff */
            {8'h00}, /* 0x7afe */
            {8'h00}, /* 0x7afd */
            {8'h00}, /* 0x7afc */
            {8'h00}, /* 0x7afb */
            {8'h00}, /* 0x7afa */
            {8'h00}, /* 0x7af9 */
            {8'h00}, /* 0x7af8 */
            {8'h00}, /* 0x7af7 */
            {8'h00}, /* 0x7af6 */
            {8'h00}, /* 0x7af5 */
            {8'h00}, /* 0x7af4 */
            {8'h00}, /* 0x7af3 */
            {8'h00}, /* 0x7af2 */
            {8'h00}, /* 0x7af1 */
            {8'h00}, /* 0x7af0 */
            {8'h00}, /* 0x7aef */
            {8'h00}, /* 0x7aee */
            {8'h00}, /* 0x7aed */
            {8'h00}, /* 0x7aec */
            {8'h00}, /* 0x7aeb */
            {8'h00}, /* 0x7aea */
            {8'h00}, /* 0x7ae9 */
            {8'h00}, /* 0x7ae8 */
            {8'h00}, /* 0x7ae7 */
            {8'h00}, /* 0x7ae6 */
            {8'h00}, /* 0x7ae5 */
            {8'h00}, /* 0x7ae4 */
            {8'h00}, /* 0x7ae3 */
            {8'h00}, /* 0x7ae2 */
            {8'h00}, /* 0x7ae1 */
            {8'h00}, /* 0x7ae0 */
            {8'h00}, /* 0x7adf */
            {8'h00}, /* 0x7ade */
            {8'h00}, /* 0x7add */
            {8'h00}, /* 0x7adc */
            {8'h00}, /* 0x7adb */
            {8'h00}, /* 0x7ada */
            {8'h00}, /* 0x7ad9 */
            {8'h00}, /* 0x7ad8 */
            {8'h00}, /* 0x7ad7 */
            {8'h00}, /* 0x7ad6 */
            {8'h00}, /* 0x7ad5 */
            {8'h00}, /* 0x7ad4 */
            {8'h00}, /* 0x7ad3 */
            {8'h00}, /* 0x7ad2 */
            {8'h00}, /* 0x7ad1 */
            {8'h00}, /* 0x7ad0 */
            {8'h00}, /* 0x7acf */
            {8'h00}, /* 0x7ace */
            {8'h00}, /* 0x7acd */
            {8'h00}, /* 0x7acc */
            {8'h00}, /* 0x7acb */
            {8'h00}, /* 0x7aca */
            {8'h00}, /* 0x7ac9 */
            {8'h00}, /* 0x7ac8 */
            {8'h00}, /* 0x7ac7 */
            {8'h00}, /* 0x7ac6 */
            {8'h00}, /* 0x7ac5 */
            {8'h00}, /* 0x7ac4 */
            {8'h00}, /* 0x7ac3 */
            {8'h00}, /* 0x7ac2 */
            {8'h00}, /* 0x7ac1 */
            {8'h00}, /* 0x7ac0 */
            {8'h00}, /* 0x7abf */
            {8'h00}, /* 0x7abe */
            {8'h00}, /* 0x7abd */
            {8'h00}, /* 0x7abc */
            {8'h00}, /* 0x7abb */
            {8'h00}, /* 0x7aba */
            {8'h00}, /* 0x7ab9 */
            {8'h00}, /* 0x7ab8 */
            {8'h00}, /* 0x7ab7 */
            {8'h00}, /* 0x7ab6 */
            {8'h00}, /* 0x7ab5 */
            {8'h00}, /* 0x7ab4 */
            {8'h00}, /* 0x7ab3 */
            {8'h00}, /* 0x7ab2 */
            {8'h00}, /* 0x7ab1 */
            {8'h00}, /* 0x7ab0 */
            {8'h00}, /* 0x7aaf */
            {8'h00}, /* 0x7aae */
            {8'h00}, /* 0x7aad */
            {8'h00}, /* 0x7aac */
            {8'h00}, /* 0x7aab */
            {8'h00}, /* 0x7aaa */
            {8'h00}, /* 0x7aa9 */
            {8'h00}, /* 0x7aa8 */
            {8'h00}, /* 0x7aa7 */
            {8'h00}, /* 0x7aa6 */
            {8'h00}, /* 0x7aa5 */
            {8'h00}, /* 0x7aa4 */
            {8'h00}, /* 0x7aa3 */
            {8'h00}, /* 0x7aa2 */
            {8'h00}, /* 0x7aa1 */
            {8'h00}, /* 0x7aa0 */
            {8'h00}, /* 0x7a9f */
            {8'h00}, /* 0x7a9e */
            {8'h00}, /* 0x7a9d */
            {8'h00}, /* 0x7a9c */
            {8'h00}, /* 0x7a9b */
            {8'h00}, /* 0x7a9a */
            {8'h00}, /* 0x7a99 */
            {8'h00}, /* 0x7a98 */
            {8'h00}, /* 0x7a97 */
            {8'h00}, /* 0x7a96 */
            {8'h00}, /* 0x7a95 */
            {8'h00}, /* 0x7a94 */
            {8'h00}, /* 0x7a93 */
            {8'h00}, /* 0x7a92 */
            {8'h00}, /* 0x7a91 */
            {8'h00}, /* 0x7a90 */
            {8'h00}, /* 0x7a8f */
            {8'h00}, /* 0x7a8e */
            {8'h00}, /* 0x7a8d */
            {8'h00}, /* 0x7a8c */
            {8'h00}, /* 0x7a8b */
            {8'h00}, /* 0x7a8a */
            {8'h00}, /* 0x7a89 */
            {8'h00}, /* 0x7a88 */
            {8'h00}, /* 0x7a87 */
            {8'h00}, /* 0x7a86 */
            {8'h00}, /* 0x7a85 */
            {8'h00}, /* 0x7a84 */
            {8'h00}, /* 0x7a83 */
            {8'h00}, /* 0x7a82 */
            {8'h00}, /* 0x7a81 */
            {8'h00}, /* 0x7a80 */
            {8'h00}, /* 0x7a7f */
            {8'h00}, /* 0x7a7e */
            {8'h00}, /* 0x7a7d */
            {8'h00}, /* 0x7a7c */
            {8'h00}, /* 0x7a7b */
            {8'h00}, /* 0x7a7a */
            {8'h00}, /* 0x7a79 */
            {8'h00}, /* 0x7a78 */
            {8'h00}, /* 0x7a77 */
            {8'h00}, /* 0x7a76 */
            {8'h00}, /* 0x7a75 */
            {8'h00}, /* 0x7a74 */
            {8'h00}, /* 0x7a73 */
            {8'h00}, /* 0x7a72 */
            {8'h00}, /* 0x7a71 */
            {8'h00}, /* 0x7a70 */
            {8'h00}, /* 0x7a6f */
            {8'h00}, /* 0x7a6e */
            {8'h00}, /* 0x7a6d */
            {8'h00}, /* 0x7a6c */
            {8'h00}, /* 0x7a6b */
            {8'h00}, /* 0x7a6a */
            {8'h00}, /* 0x7a69 */
            {8'h00}, /* 0x7a68 */
            {8'h00}, /* 0x7a67 */
            {8'h00}, /* 0x7a66 */
            {8'h00}, /* 0x7a65 */
            {8'h00}, /* 0x7a64 */
            {8'h00}, /* 0x7a63 */
            {8'h00}, /* 0x7a62 */
            {8'h00}, /* 0x7a61 */
            {8'h00}, /* 0x7a60 */
            {8'h00}, /* 0x7a5f */
            {8'h00}, /* 0x7a5e */
            {8'h00}, /* 0x7a5d */
            {8'h00}, /* 0x7a5c */
            {8'h00}, /* 0x7a5b */
            {8'h00}, /* 0x7a5a */
            {8'h00}, /* 0x7a59 */
            {8'h00}, /* 0x7a58 */
            {8'h00}, /* 0x7a57 */
            {8'h00}, /* 0x7a56 */
            {8'h00}, /* 0x7a55 */
            {8'h00}, /* 0x7a54 */
            {8'h00}, /* 0x7a53 */
            {8'h00}, /* 0x7a52 */
            {8'h00}, /* 0x7a51 */
            {8'h00}, /* 0x7a50 */
            {8'h00}, /* 0x7a4f */
            {8'h00}, /* 0x7a4e */
            {8'h00}, /* 0x7a4d */
            {8'h00}, /* 0x7a4c */
            {8'h00}, /* 0x7a4b */
            {8'h00}, /* 0x7a4a */
            {8'h00}, /* 0x7a49 */
            {8'h00}, /* 0x7a48 */
            {8'h00}, /* 0x7a47 */
            {8'h00}, /* 0x7a46 */
            {8'h00}, /* 0x7a45 */
            {8'h00}, /* 0x7a44 */
            {8'h00}, /* 0x7a43 */
            {8'h00}, /* 0x7a42 */
            {8'h00}, /* 0x7a41 */
            {8'h00}, /* 0x7a40 */
            {8'h00}, /* 0x7a3f */
            {8'h00}, /* 0x7a3e */
            {8'h00}, /* 0x7a3d */
            {8'h00}, /* 0x7a3c */
            {8'h00}, /* 0x7a3b */
            {8'h00}, /* 0x7a3a */
            {8'h00}, /* 0x7a39 */
            {8'h00}, /* 0x7a38 */
            {8'h00}, /* 0x7a37 */
            {8'h00}, /* 0x7a36 */
            {8'h00}, /* 0x7a35 */
            {8'h00}, /* 0x7a34 */
            {8'h00}, /* 0x7a33 */
            {8'h00}, /* 0x7a32 */
            {8'h00}, /* 0x7a31 */
            {8'h00}, /* 0x7a30 */
            {8'h00}, /* 0x7a2f */
            {8'h00}, /* 0x7a2e */
            {8'h00}, /* 0x7a2d */
            {8'h00}, /* 0x7a2c */
            {8'h00}, /* 0x7a2b */
            {8'h00}, /* 0x7a2a */
            {8'h00}, /* 0x7a29 */
            {8'h00}, /* 0x7a28 */
            {8'h00}, /* 0x7a27 */
            {8'h00}, /* 0x7a26 */
            {8'h00}, /* 0x7a25 */
            {8'h00}, /* 0x7a24 */
            {8'h00}, /* 0x7a23 */
            {8'h00}, /* 0x7a22 */
            {8'h00}, /* 0x7a21 */
            {8'h00}, /* 0x7a20 */
            {8'h00}, /* 0x7a1f */
            {8'h00}, /* 0x7a1e */
            {8'h00}, /* 0x7a1d */
            {8'h00}, /* 0x7a1c */
            {8'h00}, /* 0x7a1b */
            {8'h00}, /* 0x7a1a */
            {8'h00}, /* 0x7a19 */
            {8'h00}, /* 0x7a18 */
            {8'h00}, /* 0x7a17 */
            {8'h00}, /* 0x7a16 */
            {8'h00}, /* 0x7a15 */
            {8'h00}, /* 0x7a14 */
            {8'h00}, /* 0x7a13 */
            {8'h00}, /* 0x7a12 */
            {8'h00}, /* 0x7a11 */
            {8'h00}, /* 0x7a10 */
            {8'h00}, /* 0x7a0f */
            {8'h00}, /* 0x7a0e */
            {8'h00}, /* 0x7a0d */
            {8'h00}, /* 0x7a0c */
            {8'h00}, /* 0x7a0b */
            {8'h00}, /* 0x7a0a */
            {8'h00}, /* 0x7a09 */
            {8'h00}, /* 0x7a08 */
            {8'h00}, /* 0x7a07 */
            {8'h00}, /* 0x7a06 */
            {8'h00}, /* 0x7a05 */
            {8'h00}, /* 0x7a04 */
            {8'h00}, /* 0x7a03 */
            {8'h00}, /* 0x7a02 */
            {8'h00}, /* 0x7a01 */
            {8'h00}, /* 0x7a00 */
            {8'h00}, /* 0x79ff */
            {8'h00}, /* 0x79fe */
            {8'h00}, /* 0x79fd */
            {8'h00}, /* 0x79fc */
            {8'h00}, /* 0x79fb */
            {8'h00}, /* 0x79fa */
            {8'h00}, /* 0x79f9 */
            {8'h00}, /* 0x79f8 */
            {8'h00}, /* 0x79f7 */
            {8'h00}, /* 0x79f6 */
            {8'h00}, /* 0x79f5 */
            {8'h00}, /* 0x79f4 */
            {8'h00}, /* 0x79f3 */
            {8'h00}, /* 0x79f2 */
            {8'h00}, /* 0x79f1 */
            {8'h00}, /* 0x79f0 */
            {8'h00}, /* 0x79ef */
            {8'h00}, /* 0x79ee */
            {8'h00}, /* 0x79ed */
            {8'h00}, /* 0x79ec */
            {8'h00}, /* 0x79eb */
            {8'h00}, /* 0x79ea */
            {8'h00}, /* 0x79e9 */
            {8'h00}, /* 0x79e8 */
            {8'h00}, /* 0x79e7 */
            {8'h00}, /* 0x79e6 */
            {8'h00}, /* 0x79e5 */
            {8'h00}, /* 0x79e4 */
            {8'h00}, /* 0x79e3 */
            {8'h00}, /* 0x79e2 */
            {8'h00}, /* 0x79e1 */
            {8'h00}, /* 0x79e0 */
            {8'h00}, /* 0x79df */
            {8'h00}, /* 0x79de */
            {8'h00}, /* 0x79dd */
            {8'h00}, /* 0x79dc */
            {8'h00}, /* 0x79db */
            {8'h00}, /* 0x79da */
            {8'h00}, /* 0x79d9 */
            {8'h00}, /* 0x79d8 */
            {8'h00}, /* 0x79d7 */
            {8'h00}, /* 0x79d6 */
            {8'h00}, /* 0x79d5 */
            {8'h00}, /* 0x79d4 */
            {8'h00}, /* 0x79d3 */
            {8'h00}, /* 0x79d2 */
            {8'h00}, /* 0x79d1 */
            {8'h00}, /* 0x79d0 */
            {8'h00}, /* 0x79cf */
            {8'h00}, /* 0x79ce */
            {8'h00}, /* 0x79cd */
            {8'h00}, /* 0x79cc */
            {8'h00}, /* 0x79cb */
            {8'h00}, /* 0x79ca */
            {8'h00}, /* 0x79c9 */
            {8'h00}, /* 0x79c8 */
            {8'h00}, /* 0x79c7 */
            {8'h00}, /* 0x79c6 */
            {8'h00}, /* 0x79c5 */
            {8'h00}, /* 0x79c4 */
            {8'h00}, /* 0x79c3 */
            {8'h00}, /* 0x79c2 */
            {8'h00}, /* 0x79c1 */
            {8'h00}, /* 0x79c0 */
            {8'h00}, /* 0x79bf */
            {8'h00}, /* 0x79be */
            {8'h00}, /* 0x79bd */
            {8'h00}, /* 0x79bc */
            {8'h00}, /* 0x79bb */
            {8'h00}, /* 0x79ba */
            {8'h00}, /* 0x79b9 */
            {8'h00}, /* 0x79b8 */
            {8'h00}, /* 0x79b7 */
            {8'h00}, /* 0x79b6 */
            {8'h00}, /* 0x79b5 */
            {8'h00}, /* 0x79b4 */
            {8'h00}, /* 0x79b3 */
            {8'h00}, /* 0x79b2 */
            {8'h00}, /* 0x79b1 */
            {8'h00}, /* 0x79b0 */
            {8'h00}, /* 0x79af */
            {8'h00}, /* 0x79ae */
            {8'h00}, /* 0x79ad */
            {8'h00}, /* 0x79ac */
            {8'h00}, /* 0x79ab */
            {8'h00}, /* 0x79aa */
            {8'h00}, /* 0x79a9 */
            {8'h00}, /* 0x79a8 */
            {8'h00}, /* 0x79a7 */
            {8'h00}, /* 0x79a6 */
            {8'h00}, /* 0x79a5 */
            {8'h00}, /* 0x79a4 */
            {8'h00}, /* 0x79a3 */
            {8'h00}, /* 0x79a2 */
            {8'h00}, /* 0x79a1 */
            {8'h00}, /* 0x79a0 */
            {8'h00}, /* 0x799f */
            {8'h00}, /* 0x799e */
            {8'h00}, /* 0x799d */
            {8'h00}, /* 0x799c */
            {8'h00}, /* 0x799b */
            {8'h00}, /* 0x799a */
            {8'h00}, /* 0x7999 */
            {8'h00}, /* 0x7998 */
            {8'h00}, /* 0x7997 */
            {8'h00}, /* 0x7996 */
            {8'h00}, /* 0x7995 */
            {8'h00}, /* 0x7994 */
            {8'h00}, /* 0x7993 */
            {8'h00}, /* 0x7992 */
            {8'h00}, /* 0x7991 */
            {8'h00}, /* 0x7990 */
            {8'h00}, /* 0x798f */
            {8'h00}, /* 0x798e */
            {8'h00}, /* 0x798d */
            {8'h00}, /* 0x798c */
            {8'h00}, /* 0x798b */
            {8'h00}, /* 0x798a */
            {8'h00}, /* 0x7989 */
            {8'h00}, /* 0x7988 */
            {8'h00}, /* 0x7987 */
            {8'h00}, /* 0x7986 */
            {8'h00}, /* 0x7985 */
            {8'h00}, /* 0x7984 */
            {8'h00}, /* 0x7983 */
            {8'h00}, /* 0x7982 */
            {8'h00}, /* 0x7981 */
            {8'h00}, /* 0x7980 */
            {8'h00}, /* 0x797f */
            {8'h00}, /* 0x797e */
            {8'h00}, /* 0x797d */
            {8'h00}, /* 0x797c */
            {8'h00}, /* 0x797b */
            {8'h00}, /* 0x797a */
            {8'h00}, /* 0x7979 */
            {8'h00}, /* 0x7978 */
            {8'h00}, /* 0x7977 */
            {8'h00}, /* 0x7976 */
            {8'h00}, /* 0x7975 */
            {8'h00}, /* 0x7974 */
            {8'h00}, /* 0x7973 */
            {8'h00}, /* 0x7972 */
            {8'h00}, /* 0x7971 */
            {8'h00}, /* 0x7970 */
            {8'h00}, /* 0x796f */
            {8'h00}, /* 0x796e */
            {8'h00}, /* 0x796d */
            {8'h00}, /* 0x796c */
            {8'h00}, /* 0x796b */
            {8'h00}, /* 0x796a */
            {8'h00}, /* 0x7969 */
            {8'h00}, /* 0x7968 */
            {8'h00}, /* 0x7967 */
            {8'h00}, /* 0x7966 */
            {8'h00}, /* 0x7965 */
            {8'h00}, /* 0x7964 */
            {8'h00}, /* 0x7963 */
            {8'h00}, /* 0x7962 */
            {8'h00}, /* 0x7961 */
            {8'h00}, /* 0x7960 */
            {8'h00}, /* 0x795f */
            {8'h00}, /* 0x795e */
            {8'h00}, /* 0x795d */
            {8'h00}, /* 0x795c */
            {8'h00}, /* 0x795b */
            {8'h00}, /* 0x795a */
            {8'h00}, /* 0x7959 */
            {8'h00}, /* 0x7958 */
            {8'h00}, /* 0x7957 */
            {8'h00}, /* 0x7956 */
            {8'h00}, /* 0x7955 */
            {8'h00}, /* 0x7954 */
            {8'h00}, /* 0x7953 */
            {8'h00}, /* 0x7952 */
            {8'h00}, /* 0x7951 */
            {8'h00}, /* 0x7950 */
            {8'h00}, /* 0x794f */
            {8'h00}, /* 0x794e */
            {8'h00}, /* 0x794d */
            {8'h00}, /* 0x794c */
            {8'h00}, /* 0x794b */
            {8'h00}, /* 0x794a */
            {8'h00}, /* 0x7949 */
            {8'h00}, /* 0x7948 */
            {8'h00}, /* 0x7947 */
            {8'h00}, /* 0x7946 */
            {8'h00}, /* 0x7945 */
            {8'h00}, /* 0x7944 */
            {8'h00}, /* 0x7943 */
            {8'h00}, /* 0x7942 */
            {8'h00}, /* 0x7941 */
            {8'h00}, /* 0x7940 */
            {8'h00}, /* 0x793f */
            {8'h00}, /* 0x793e */
            {8'h00}, /* 0x793d */
            {8'h00}, /* 0x793c */
            {8'h00}, /* 0x793b */
            {8'h00}, /* 0x793a */
            {8'h00}, /* 0x7939 */
            {8'h00}, /* 0x7938 */
            {8'h00}, /* 0x7937 */
            {8'h00}, /* 0x7936 */
            {8'h00}, /* 0x7935 */
            {8'h00}, /* 0x7934 */
            {8'h00}, /* 0x7933 */
            {8'h00}, /* 0x7932 */
            {8'h00}, /* 0x7931 */
            {8'h00}, /* 0x7930 */
            {8'h00}, /* 0x792f */
            {8'h00}, /* 0x792e */
            {8'h00}, /* 0x792d */
            {8'h00}, /* 0x792c */
            {8'h00}, /* 0x792b */
            {8'h00}, /* 0x792a */
            {8'h00}, /* 0x7929 */
            {8'h00}, /* 0x7928 */
            {8'h00}, /* 0x7927 */
            {8'h00}, /* 0x7926 */
            {8'h00}, /* 0x7925 */
            {8'h00}, /* 0x7924 */
            {8'h00}, /* 0x7923 */
            {8'h00}, /* 0x7922 */
            {8'h00}, /* 0x7921 */
            {8'h00}, /* 0x7920 */
            {8'h00}, /* 0x791f */
            {8'h00}, /* 0x791e */
            {8'h00}, /* 0x791d */
            {8'h00}, /* 0x791c */
            {8'h00}, /* 0x791b */
            {8'h00}, /* 0x791a */
            {8'h00}, /* 0x7919 */
            {8'h00}, /* 0x7918 */
            {8'h00}, /* 0x7917 */
            {8'h00}, /* 0x7916 */
            {8'h00}, /* 0x7915 */
            {8'h00}, /* 0x7914 */
            {8'h00}, /* 0x7913 */
            {8'h00}, /* 0x7912 */
            {8'h00}, /* 0x7911 */
            {8'h00}, /* 0x7910 */
            {8'h00}, /* 0x790f */
            {8'h00}, /* 0x790e */
            {8'h00}, /* 0x790d */
            {8'h00}, /* 0x790c */
            {8'h00}, /* 0x790b */
            {8'h00}, /* 0x790a */
            {8'h00}, /* 0x7909 */
            {8'h00}, /* 0x7908 */
            {8'h00}, /* 0x7907 */
            {8'h00}, /* 0x7906 */
            {8'h00}, /* 0x7905 */
            {8'h00}, /* 0x7904 */
            {8'h00}, /* 0x7903 */
            {8'h00}, /* 0x7902 */
            {8'h00}, /* 0x7901 */
            {8'h00}, /* 0x7900 */
            {8'h00}, /* 0x78ff */
            {8'h00}, /* 0x78fe */
            {8'h00}, /* 0x78fd */
            {8'h00}, /* 0x78fc */
            {8'h00}, /* 0x78fb */
            {8'h00}, /* 0x78fa */
            {8'h00}, /* 0x78f9 */
            {8'h00}, /* 0x78f8 */
            {8'h00}, /* 0x78f7 */
            {8'h00}, /* 0x78f6 */
            {8'h00}, /* 0x78f5 */
            {8'h00}, /* 0x78f4 */
            {8'h00}, /* 0x78f3 */
            {8'h00}, /* 0x78f2 */
            {8'h00}, /* 0x78f1 */
            {8'h00}, /* 0x78f0 */
            {8'h00}, /* 0x78ef */
            {8'h00}, /* 0x78ee */
            {8'h00}, /* 0x78ed */
            {8'h00}, /* 0x78ec */
            {8'h00}, /* 0x78eb */
            {8'h00}, /* 0x78ea */
            {8'h00}, /* 0x78e9 */
            {8'h00}, /* 0x78e8 */
            {8'h00}, /* 0x78e7 */
            {8'h00}, /* 0x78e6 */
            {8'h00}, /* 0x78e5 */
            {8'h00}, /* 0x78e4 */
            {8'h00}, /* 0x78e3 */
            {8'h00}, /* 0x78e2 */
            {8'h00}, /* 0x78e1 */
            {8'h00}, /* 0x78e0 */
            {8'h00}, /* 0x78df */
            {8'h00}, /* 0x78de */
            {8'h00}, /* 0x78dd */
            {8'h00}, /* 0x78dc */
            {8'h00}, /* 0x78db */
            {8'h00}, /* 0x78da */
            {8'h00}, /* 0x78d9 */
            {8'h00}, /* 0x78d8 */
            {8'h00}, /* 0x78d7 */
            {8'h00}, /* 0x78d6 */
            {8'h00}, /* 0x78d5 */
            {8'h00}, /* 0x78d4 */
            {8'h00}, /* 0x78d3 */
            {8'h00}, /* 0x78d2 */
            {8'h00}, /* 0x78d1 */
            {8'h00}, /* 0x78d0 */
            {8'h00}, /* 0x78cf */
            {8'h00}, /* 0x78ce */
            {8'h00}, /* 0x78cd */
            {8'h00}, /* 0x78cc */
            {8'h00}, /* 0x78cb */
            {8'h00}, /* 0x78ca */
            {8'h00}, /* 0x78c9 */
            {8'h00}, /* 0x78c8 */
            {8'h00}, /* 0x78c7 */
            {8'h00}, /* 0x78c6 */
            {8'h00}, /* 0x78c5 */
            {8'h00}, /* 0x78c4 */
            {8'h00}, /* 0x78c3 */
            {8'h00}, /* 0x78c2 */
            {8'h00}, /* 0x78c1 */
            {8'h00}, /* 0x78c0 */
            {8'h00}, /* 0x78bf */
            {8'h00}, /* 0x78be */
            {8'h00}, /* 0x78bd */
            {8'h00}, /* 0x78bc */
            {8'h00}, /* 0x78bb */
            {8'h00}, /* 0x78ba */
            {8'h00}, /* 0x78b9 */
            {8'h00}, /* 0x78b8 */
            {8'h00}, /* 0x78b7 */
            {8'h00}, /* 0x78b6 */
            {8'h00}, /* 0x78b5 */
            {8'h00}, /* 0x78b4 */
            {8'h00}, /* 0x78b3 */
            {8'h00}, /* 0x78b2 */
            {8'h00}, /* 0x78b1 */
            {8'h00}, /* 0x78b0 */
            {8'h00}, /* 0x78af */
            {8'h00}, /* 0x78ae */
            {8'h00}, /* 0x78ad */
            {8'h00}, /* 0x78ac */
            {8'h00}, /* 0x78ab */
            {8'h00}, /* 0x78aa */
            {8'h00}, /* 0x78a9 */
            {8'h00}, /* 0x78a8 */
            {8'h00}, /* 0x78a7 */
            {8'h00}, /* 0x78a6 */
            {8'h00}, /* 0x78a5 */
            {8'h00}, /* 0x78a4 */
            {8'h00}, /* 0x78a3 */
            {8'h00}, /* 0x78a2 */
            {8'h00}, /* 0x78a1 */
            {8'h00}, /* 0x78a0 */
            {8'h00}, /* 0x789f */
            {8'h00}, /* 0x789e */
            {8'h00}, /* 0x789d */
            {8'h00}, /* 0x789c */
            {8'h00}, /* 0x789b */
            {8'h00}, /* 0x789a */
            {8'h00}, /* 0x7899 */
            {8'h00}, /* 0x7898 */
            {8'h00}, /* 0x7897 */
            {8'h00}, /* 0x7896 */
            {8'h00}, /* 0x7895 */
            {8'h00}, /* 0x7894 */
            {8'h00}, /* 0x7893 */
            {8'h00}, /* 0x7892 */
            {8'h00}, /* 0x7891 */
            {8'h00}, /* 0x7890 */
            {8'h00}, /* 0x788f */
            {8'h00}, /* 0x788e */
            {8'h00}, /* 0x788d */
            {8'h00}, /* 0x788c */
            {8'h00}, /* 0x788b */
            {8'h00}, /* 0x788a */
            {8'h00}, /* 0x7889 */
            {8'h00}, /* 0x7888 */
            {8'h00}, /* 0x7887 */
            {8'h00}, /* 0x7886 */
            {8'h00}, /* 0x7885 */
            {8'h00}, /* 0x7884 */
            {8'h00}, /* 0x7883 */
            {8'h00}, /* 0x7882 */
            {8'h00}, /* 0x7881 */
            {8'h00}, /* 0x7880 */
            {8'h00}, /* 0x787f */
            {8'h00}, /* 0x787e */
            {8'h00}, /* 0x787d */
            {8'h00}, /* 0x787c */
            {8'h00}, /* 0x787b */
            {8'h00}, /* 0x787a */
            {8'h00}, /* 0x7879 */
            {8'h00}, /* 0x7878 */
            {8'h00}, /* 0x7877 */
            {8'h00}, /* 0x7876 */
            {8'h00}, /* 0x7875 */
            {8'h00}, /* 0x7874 */
            {8'h00}, /* 0x7873 */
            {8'h00}, /* 0x7872 */
            {8'h00}, /* 0x7871 */
            {8'h00}, /* 0x7870 */
            {8'h00}, /* 0x786f */
            {8'h00}, /* 0x786e */
            {8'h00}, /* 0x786d */
            {8'h00}, /* 0x786c */
            {8'h00}, /* 0x786b */
            {8'h00}, /* 0x786a */
            {8'h00}, /* 0x7869 */
            {8'h00}, /* 0x7868 */
            {8'h00}, /* 0x7867 */
            {8'h00}, /* 0x7866 */
            {8'h00}, /* 0x7865 */
            {8'h00}, /* 0x7864 */
            {8'h00}, /* 0x7863 */
            {8'h00}, /* 0x7862 */
            {8'h00}, /* 0x7861 */
            {8'h00}, /* 0x7860 */
            {8'h00}, /* 0x785f */
            {8'h00}, /* 0x785e */
            {8'h00}, /* 0x785d */
            {8'h00}, /* 0x785c */
            {8'h00}, /* 0x785b */
            {8'h00}, /* 0x785a */
            {8'h00}, /* 0x7859 */
            {8'h00}, /* 0x7858 */
            {8'h00}, /* 0x7857 */
            {8'h00}, /* 0x7856 */
            {8'h00}, /* 0x7855 */
            {8'h00}, /* 0x7854 */
            {8'h00}, /* 0x7853 */
            {8'h00}, /* 0x7852 */
            {8'h00}, /* 0x7851 */
            {8'h00}, /* 0x7850 */
            {8'h00}, /* 0x784f */
            {8'h00}, /* 0x784e */
            {8'h00}, /* 0x784d */
            {8'h00}, /* 0x784c */
            {8'h00}, /* 0x784b */
            {8'h00}, /* 0x784a */
            {8'h00}, /* 0x7849 */
            {8'h00}, /* 0x7848 */
            {8'h00}, /* 0x7847 */
            {8'h00}, /* 0x7846 */
            {8'h00}, /* 0x7845 */
            {8'h00}, /* 0x7844 */
            {8'h00}, /* 0x7843 */
            {8'h00}, /* 0x7842 */
            {8'h00}, /* 0x7841 */
            {8'h00}, /* 0x7840 */
            {8'h00}, /* 0x783f */
            {8'h00}, /* 0x783e */
            {8'h00}, /* 0x783d */
            {8'h00}, /* 0x783c */
            {8'h00}, /* 0x783b */
            {8'h00}, /* 0x783a */
            {8'h00}, /* 0x7839 */
            {8'h00}, /* 0x7838 */
            {8'h00}, /* 0x7837 */
            {8'h00}, /* 0x7836 */
            {8'h00}, /* 0x7835 */
            {8'h00}, /* 0x7834 */
            {8'h00}, /* 0x7833 */
            {8'h00}, /* 0x7832 */
            {8'h00}, /* 0x7831 */
            {8'h00}, /* 0x7830 */
            {8'h00}, /* 0x782f */
            {8'h00}, /* 0x782e */
            {8'h00}, /* 0x782d */
            {8'h00}, /* 0x782c */
            {8'h00}, /* 0x782b */
            {8'h00}, /* 0x782a */
            {8'h00}, /* 0x7829 */
            {8'h00}, /* 0x7828 */
            {8'h00}, /* 0x7827 */
            {8'h00}, /* 0x7826 */
            {8'h00}, /* 0x7825 */
            {8'h00}, /* 0x7824 */
            {8'h00}, /* 0x7823 */
            {8'h00}, /* 0x7822 */
            {8'h00}, /* 0x7821 */
            {8'h00}, /* 0x7820 */
            {8'h00}, /* 0x781f */
            {8'h00}, /* 0x781e */
            {8'h00}, /* 0x781d */
            {8'h00}, /* 0x781c */
            {8'h00}, /* 0x781b */
            {8'h00}, /* 0x781a */
            {8'h00}, /* 0x7819 */
            {8'h00}, /* 0x7818 */
            {8'h00}, /* 0x7817 */
            {8'h00}, /* 0x7816 */
            {8'h00}, /* 0x7815 */
            {8'h00}, /* 0x7814 */
            {8'h00}, /* 0x7813 */
            {8'h00}, /* 0x7812 */
            {8'h00}, /* 0x7811 */
            {8'h00}, /* 0x7810 */
            {8'h00}, /* 0x780f */
            {8'h00}, /* 0x780e */
            {8'h00}, /* 0x780d */
            {8'h00}, /* 0x780c */
            {8'h00}, /* 0x780b */
            {8'h00}, /* 0x780a */
            {8'h00}, /* 0x7809 */
            {8'h00}, /* 0x7808 */
            {8'h00}, /* 0x7807 */
            {8'h00}, /* 0x7806 */
            {8'h00}, /* 0x7805 */
            {8'h00}, /* 0x7804 */
            {8'h00}, /* 0x7803 */
            {8'h00}, /* 0x7802 */
            {8'h00}, /* 0x7801 */
            {8'h00}, /* 0x7800 */
            {8'h00}, /* 0x77ff */
            {8'h00}, /* 0x77fe */
            {8'h00}, /* 0x77fd */
            {8'h00}, /* 0x77fc */
            {8'h00}, /* 0x77fb */
            {8'h00}, /* 0x77fa */
            {8'h00}, /* 0x77f9 */
            {8'h00}, /* 0x77f8 */
            {8'h00}, /* 0x77f7 */
            {8'h00}, /* 0x77f6 */
            {8'h00}, /* 0x77f5 */
            {8'h00}, /* 0x77f4 */
            {8'h00}, /* 0x77f3 */
            {8'h00}, /* 0x77f2 */
            {8'h00}, /* 0x77f1 */
            {8'h00}, /* 0x77f0 */
            {8'h00}, /* 0x77ef */
            {8'h00}, /* 0x77ee */
            {8'h00}, /* 0x77ed */
            {8'h00}, /* 0x77ec */
            {8'h00}, /* 0x77eb */
            {8'h00}, /* 0x77ea */
            {8'h00}, /* 0x77e9 */
            {8'h00}, /* 0x77e8 */
            {8'h00}, /* 0x77e7 */
            {8'h00}, /* 0x77e6 */
            {8'h00}, /* 0x77e5 */
            {8'h00}, /* 0x77e4 */
            {8'h00}, /* 0x77e3 */
            {8'h00}, /* 0x77e2 */
            {8'h00}, /* 0x77e1 */
            {8'h00}, /* 0x77e0 */
            {8'h00}, /* 0x77df */
            {8'h00}, /* 0x77de */
            {8'h00}, /* 0x77dd */
            {8'h00}, /* 0x77dc */
            {8'h00}, /* 0x77db */
            {8'h00}, /* 0x77da */
            {8'h00}, /* 0x77d9 */
            {8'h00}, /* 0x77d8 */
            {8'h00}, /* 0x77d7 */
            {8'h00}, /* 0x77d6 */
            {8'h00}, /* 0x77d5 */
            {8'h00}, /* 0x77d4 */
            {8'h00}, /* 0x77d3 */
            {8'h00}, /* 0x77d2 */
            {8'h00}, /* 0x77d1 */
            {8'h00}, /* 0x77d0 */
            {8'h00}, /* 0x77cf */
            {8'h00}, /* 0x77ce */
            {8'h00}, /* 0x77cd */
            {8'h00}, /* 0x77cc */
            {8'h00}, /* 0x77cb */
            {8'h00}, /* 0x77ca */
            {8'h00}, /* 0x77c9 */
            {8'h00}, /* 0x77c8 */
            {8'h00}, /* 0x77c7 */
            {8'h00}, /* 0x77c6 */
            {8'h00}, /* 0x77c5 */
            {8'h00}, /* 0x77c4 */
            {8'h00}, /* 0x77c3 */
            {8'h00}, /* 0x77c2 */
            {8'h00}, /* 0x77c1 */
            {8'h00}, /* 0x77c0 */
            {8'h00}, /* 0x77bf */
            {8'h00}, /* 0x77be */
            {8'h00}, /* 0x77bd */
            {8'h00}, /* 0x77bc */
            {8'h00}, /* 0x77bb */
            {8'h00}, /* 0x77ba */
            {8'h00}, /* 0x77b9 */
            {8'h00}, /* 0x77b8 */
            {8'h00}, /* 0x77b7 */
            {8'h00}, /* 0x77b6 */
            {8'h00}, /* 0x77b5 */
            {8'h00}, /* 0x77b4 */
            {8'h00}, /* 0x77b3 */
            {8'h00}, /* 0x77b2 */
            {8'h00}, /* 0x77b1 */
            {8'h00}, /* 0x77b0 */
            {8'h00}, /* 0x77af */
            {8'h00}, /* 0x77ae */
            {8'h00}, /* 0x77ad */
            {8'h00}, /* 0x77ac */
            {8'h00}, /* 0x77ab */
            {8'h00}, /* 0x77aa */
            {8'h00}, /* 0x77a9 */
            {8'h00}, /* 0x77a8 */
            {8'h00}, /* 0x77a7 */
            {8'h00}, /* 0x77a6 */
            {8'h00}, /* 0x77a5 */
            {8'h00}, /* 0x77a4 */
            {8'h00}, /* 0x77a3 */
            {8'h00}, /* 0x77a2 */
            {8'h00}, /* 0x77a1 */
            {8'h00}, /* 0x77a0 */
            {8'h00}, /* 0x779f */
            {8'h00}, /* 0x779e */
            {8'h00}, /* 0x779d */
            {8'h00}, /* 0x779c */
            {8'h00}, /* 0x779b */
            {8'h00}, /* 0x779a */
            {8'h00}, /* 0x7799 */
            {8'h00}, /* 0x7798 */
            {8'h00}, /* 0x7797 */
            {8'h00}, /* 0x7796 */
            {8'h00}, /* 0x7795 */
            {8'h00}, /* 0x7794 */
            {8'h00}, /* 0x7793 */
            {8'h00}, /* 0x7792 */
            {8'h00}, /* 0x7791 */
            {8'h00}, /* 0x7790 */
            {8'h00}, /* 0x778f */
            {8'h00}, /* 0x778e */
            {8'h00}, /* 0x778d */
            {8'h00}, /* 0x778c */
            {8'h00}, /* 0x778b */
            {8'h00}, /* 0x778a */
            {8'h00}, /* 0x7789 */
            {8'h00}, /* 0x7788 */
            {8'h00}, /* 0x7787 */
            {8'h00}, /* 0x7786 */
            {8'h00}, /* 0x7785 */
            {8'h00}, /* 0x7784 */
            {8'h00}, /* 0x7783 */
            {8'h00}, /* 0x7782 */
            {8'h00}, /* 0x7781 */
            {8'h00}, /* 0x7780 */
            {8'h00}, /* 0x777f */
            {8'h00}, /* 0x777e */
            {8'h00}, /* 0x777d */
            {8'h00}, /* 0x777c */
            {8'h00}, /* 0x777b */
            {8'h00}, /* 0x777a */
            {8'h00}, /* 0x7779 */
            {8'h00}, /* 0x7778 */
            {8'h00}, /* 0x7777 */
            {8'h00}, /* 0x7776 */
            {8'h00}, /* 0x7775 */
            {8'h00}, /* 0x7774 */
            {8'h00}, /* 0x7773 */
            {8'h00}, /* 0x7772 */
            {8'h00}, /* 0x7771 */
            {8'h00}, /* 0x7770 */
            {8'h00}, /* 0x776f */
            {8'h00}, /* 0x776e */
            {8'h00}, /* 0x776d */
            {8'h00}, /* 0x776c */
            {8'h00}, /* 0x776b */
            {8'h00}, /* 0x776a */
            {8'h00}, /* 0x7769 */
            {8'h00}, /* 0x7768 */
            {8'h00}, /* 0x7767 */
            {8'h00}, /* 0x7766 */
            {8'h00}, /* 0x7765 */
            {8'h00}, /* 0x7764 */
            {8'h00}, /* 0x7763 */
            {8'h00}, /* 0x7762 */
            {8'h00}, /* 0x7761 */
            {8'h00}, /* 0x7760 */
            {8'h00}, /* 0x775f */
            {8'h00}, /* 0x775e */
            {8'h00}, /* 0x775d */
            {8'h00}, /* 0x775c */
            {8'h00}, /* 0x775b */
            {8'h00}, /* 0x775a */
            {8'h00}, /* 0x7759 */
            {8'h00}, /* 0x7758 */
            {8'h00}, /* 0x7757 */
            {8'h00}, /* 0x7756 */
            {8'h00}, /* 0x7755 */
            {8'h00}, /* 0x7754 */
            {8'h00}, /* 0x7753 */
            {8'h00}, /* 0x7752 */
            {8'h00}, /* 0x7751 */
            {8'h00}, /* 0x7750 */
            {8'h00}, /* 0x774f */
            {8'h00}, /* 0x774e */
            {8'h00}, /* 0x774d */
            {8'h00}, /* 0x774c */
            {8'h00}, /* 0x774b */
            {8'h00}, /* 0x774a */
            {8'h00}, /* 0x7749 */
            {8'h00}, /* 0x7748 */
            {8'h00}, /* 0x7747 */
            {8'h00}, /* 0x7746 */
            {8'h00}, /* 0x7745 */
            {8'h00}, /* 0x7744 */
            {8'h00}, /* 0x7743 */
            {8'h00}, /* 0x7742 */
            {8'h00}, /* 0x7741 */
            {8'h00}, /* 0x7740 */
            {8'h00}, /* 0x773f */
            {8'h00}, /* 0x773e */
            {8'h00}, /* 0x773d */
            {8'h00}, /* 0x773c */
            {8'h00}, /* 0x773b */
            {8'h00}, /* 0x773a */
            {8'h00}, /* 0x7739 */
            {8'h00}, /* 0x7738 */
            {8'h00}, /* 0x7737 */
            {8'h00}, /* 0x7736 */
            {8'h00}, /* 0x7735 */
            {8'h00}, /* 0x7734 */
            {8'h00}, /* 0x7733 */
            {8'h00}, /* 0x7732 */
            {8'h00}, /* 0x7731 */
            {8'h00}, /* 0x7730 */
            {8'h00}, /* 0x772f */
            {8'h00}, /* 0x772e */
            {8'h00}, /* 0x772d */
            {8'h00}, /* 0x772c */
            {8'h00}, /* 0x772b */
            {8'h00}, /* 0x772a */
            {8'h00}, /* 0x7729 */
            {8'h00}, /* 0x7728 */
            {8'h00}, /* 0x7727 */
            {8'h00}, /* 0x7726 */
            {8'h00}, /* 0x7725 */
            {8'h00}, /* 0x7724 */
            {8'h00}, /* 0x7723 */
            {8'h00}, /* 0x7722 */
            {8'h00}, /* 0x7721 */
            {8'h00}, /* 0x7720 */
            {8'h00}, /* 0x771f */
            {8'h00}, /* 0x771e */
            {8'h00}, /* 0x771d */
            {8'h00}, /* 0x771c */
            {8'h00}, /* 0x771b */
            {8'h00}, /* 0x771a */
            {8'h00}, /* 0x7719 */
            {8'h00}, /* 0x7718 */
            {8'h00}, /* 0x7717 */
            {8'h00}, /* 0x7716 */
            {8'h00}, /* 0x7715 */
            {8'h00}, /* 0x7714 */
            {8'h00}, /* 0x7713 */
            {8'h00}, /* 0x7712 */
            {8'h00}, /* 0x7711 */
            {8'h00}, /* 0x7710 */
            {8'h00}, /* 0x770f */
            {8'h00}, /* 0x770e */
            {8'h00}, /* 0x770d */
            {8'h00}, /* 0x770c */
            {8'h00}, /* 0x770b */
            {8'h00}, /* 0x770a */
            {8'h00}, /* 0x7709 */
            {8'h00}, /* 0x7708 */
            {8'h00}, /* 0x7707 */
            {8'h00}, /* 0x7706 */
            {8'h00}, /* 0x7705 */
            {8'h00}, /* 0x7704 */
            {8'h00}, /* 0x7703 */
            {8'h00}, /* 0x7702 */
            {8'h00}, /* 0x7701 */
            {8'h00}, /* 0x7700 */
            {8'h00}, /* 0x76ff */
            {8'h00}, /* 0x76fe */
            {8'h00}, /* 0x76fd */
            {8'h00}, /* 0x76fc */
            {8'h00}, /* 0x76fb */
            {8'h00}, /* 0x76fa */
            {8'h00}, /* 0x76f9 */
            {8'h00}, /* 0x76f8 */
            {8'h00}, /* 0x76f7 */
            {8'h00}, /* 0x76f6 */
            {8'h00}, /* 0x76f5 */
            {8'h00}, /* 0x76f4 */
            {8'h00}, /* 0x76f3 */
            {8'h00}, /* 0x76f2 */
            {8'h00}, /* 0x76f1 */
            {8'h00}, /* 0x76f0 */
            {8'h00}, /* 0x76ef */
            {8'h00}, /* 0x76ee */
            {8'h00}, /* 0x76ed */
            {8'h00}, /* 0x76ec */
            {8'h00}, /* 0x76eb */
            {8'h00}, /* 0x76ea */
            {8'h00}, /* 0x76e9 */
            {8'h00}, /* 0x76e8 */
            {8'h00}, /* 0x76e7 */
            {8'h00}, /* 0x76e6 */
            {8'h00}, /* 0x76e5 */
            {8'h00}, /* 0x76e4 */
            {8'h00}, /* 0x76e3 */
            {8'h00}, /* 0x76e2 */
            {8'h00}, /* 0x76e1 */
            {8'h00}, /* 0x76e0 */
            {8'h00}, /* 0x76df */
            {8'h00}, /* 0x76de */
            {8'h00}, /* 0x76dd */
            {8'h00}, /* 0x76dc */
            {8'h00}, /* 0x76db */
            {8'h00}, /* 0x76da */
            {8'h00}, /* 0x76d9 */
            {8'h00}, /* 0x76d8 */
            {8'h00}, /* 0x76d7 */
            {8'h00}, /* 0x76d6 */
            {8'h00}, /* 0x76d5 */
            {8'h00}, /* 0x76d4 */
            {8'h00}, /* 0x76d3 */
            {8'h00}, /* 0x76d2 */
            {8'h00}, /* 0x76d1 */
            {8'h00}, /* 0x76d0 */
            {8'h00}, /* 0x76cf */
            {8'h00}, /* 0x76ce */
            {8'h00}, /* 0x76cd */
            {8'h00}, /* 0x76cc */
            {8'h00}, /* 0x76cb */
            {8'h00}, /* 0x76ca */
            {8'h00}, /* 0x76c9 */
            {8'h00}, /* 0x76c8 */
            {8'h00}, /* 0x76c7 */
            {8'h00}, /* 0x76c6 */
            {8'h00}, /* 0x76c5 */
            {8'h00}, /* 0x76c4 */
            {8'h00}, /* 0x76c3 */
            {8'h00}, /* 0x76c2 */
            {8'h00}, /* 0x76c1 */
            {8'h00}, /* 0x76c0 */
            {8'h00}, /* 0x76bf */
            {8'h00}, /* 0x76be */
            {8'h00}, /* 0x76bd */
            {8'h00}, /* 0x76bc */
            {8'h00}, /* 0x76bb */
            {8'h00}, /* 0x76ba */
            {8'h00}, /* 0x76b9 */
            {8'h00}, /* 0x76b8 */
            {8'h00}, /* 0x76b7 */
            {8'h00}, /* 0x76b6 */
            {8'h00}, /* 0x76b5 */
            {8'h00}, /* 0x76b4 */
            {8'h00}, /* 0x76b3 */
            {8'h00}, /* 0x76b2 */
            {8'h00}, /* 0x76b1 */
            {8'h00}, /* 0x76b0 */
            {8'h00}, /* 0x76af */
            {8'h00}, /* 0x76ae */
            {8'h00}, /* 0x76ad */
            {8'h00}, /* 0x76ac */
            {8'h00}, /* 0x76ab */
            {8'h00}, /* 0x76aa */
            {8'h00}, /* 0x76a9 */
            {8'h00}, /* 0x76a8 */
            {8'h00}, /* 0x76a7 */
            {8'h00}, /* 0x76a6 */
            {8'h00}, /* 0x76a5 */
            {8'h00}, /* 0x76a4 */
            {8'h00}, /* 0x76a3 */
            {8'h00}, /* 0x76a2 */
            {8'h00}, /* 0x76a1 */
            {8'h00}, /* 0x76a0 */
            {8'h00}, /* 0x769f */
            {8'h00}, /* 0x769e */
            {8'h00}, /* 0x769d */
            {8'h00}, /* 0x769c */
            {8'h00}, /* 0x769b */
            {8'h00}, /* 0x769a */
            {8'h00}, /* 0x7699 */
            {8'h00}, /* 0x7698 */
            {8'h00}, /* 0x7697 */
            {8'h00}, /* 0x7696 */
            {8'h00}, /* 0x7695 */
            {8'h00}, /* 0x7694 */
            {8'h00}, /* 0x7693 */
            {8'h00}, /* 0x7692 */
            {8'h00}, /* 0x7691 */
            {8'h00}, /* 0x7690 */
            {8'h00}, /* 0x768f */
            {8'h00}, /* 0x768e */
            {8'h00}, /* 0x768d */
            {8'h00}, /* 0x768c */
            {8'h00}, /* 0x768b */
            {8'h00}, /* 0x768a */
            {8'h00}, /* 0x7689 */
            {8'h00}, /* 0x7688 */
            {8'h00}, /* 0x7687 */
            {8'h00}, /* 0x7686 */
            {8'h00}, /* 0x7685 */
            {8'h00}, /* 0x7684 */
            {8'h00}, /* 0x7683 */
            {8'h00}, /* 0x7682 */
            {8'h00}, /* 0x7681 */
            {8'h00}, /* 0x7680 */
            {8'h00}, /* 0x767f */
            {8'h00}, /* 0x767e */
            {8'h00}, /* 0x767d */
            {8'h00}, /* 0x767c */
            {8'h00}, /* 0x767b */
            {8'h00}, /* 0x767a */
            {8'h00}, /* 0x7679 */
            {8'h00}, /* 0x7678 */
            {8'h00}, /* 0x7677 */
            {8'h00}, /* 0x7676 */
            {8'h00}, /* 0x7675 */
            {8'h00}, /* 0x7674 */
            {8'h00}, /* 0x7673 */
            {8'h00}, /* 0x7672 */
            {8'h00}, /* 0x7671 */
            {8'h00}, /* 0x7670 */
            {8'h00}, /* 0x766f */
            {8'h00}, /* 0x766e */
            {8'h00}, /* 0x766d */
            {8'h00}, /* 0x766c */
            {8'h00}, /* 0x766b */
            {8'h00}, /* 0x766a */
            {8'h00}, /* 0x7669 */
            {8'h00}, /* 0x7668 */
            {8'h00}, /* 0x7667 */
            {8'h00}, /* 0x7666 */
            {8'h00}, /* 0x7665 */
            {8'h00}, /* 0x7664 */
            {8'h00}, /* 0x7663 */
            {8'h00}, /* 0x7662 */
            {8'h00}, /* 0x7661 */
            {8'h00}, /* 0x7660 */
            {8'h00}, /* 0x765f */
            {8'h00}, /* 0x765e */
            {8'h00}, /* 0x765d */
            {8'h00}, /* 0x765c */
            {8'h00}, /* 0x765b */
            {8'h00}, /* 0x765a */
            {8'h00}, /* 0x7659 */
            {8'h00}, /* 0x7658 */
            {8'h00}, /* 0x7657 */
            {8'h00}, /* 0x7656 */
            {8'h00}, /* 0x7655 */
            {8'h00}, /* 0x7654 */
            {8'h00}, /* 0x7653 */
            {8'h00}, /* 0x7652 */
            {8'h00}, /* 0x7651 */
            {8'h00}, /* 0x7650 */
            {8'h00}, /* 0x764f */
            {8'h00}, /* 0x764e */
            {8'h00}, /* 0x764d */
            {8'h00}, /* 0x764c */
            {8'h00}, /* 0x764b */
            {8'h00}, /* 0x764a */
            {8'h00}, /* 0x7649 */
            {8'h00}, /* 0x7648 */
            {8'h00}, /* 0x7647 */
            {8'h00}, /* 0x7646 */
            {8'h00}, /* 0x7645 */
            {8'h00}, /* 0x7644 */
            {8'h00}, /* 0x7643 */
            {8'h00}, /* 0x7642 */
            {8'h00}, /* 0x7641 */
            {8'h00}, /* 0x7640 */
            {8'h00}, /* 0x763f */
            {8'h00}, /* 0x763e */
            {8'h00}, /* 0x763d */
            {8'h00}, /* 0x763c */
            {8'h00}, /* 0x763b */
            {8'h00}, /* 0x763a */
            {8'h00}, /* 0x7639 */
            {8'h00}, /* 0x7638 */
            {8'h00}, /* 0x7637 */
            {8'h00}, /* 0x7636 */
            {8'h00}, /* 0x7635 */
            {8'h00}, /* 0x7634 */
            {8'h00}, /* 0x7633 */
            {8'h00}, /* 0x7632 */
            {8'h00}, /* 0x7631 */
            {8'h00}, /* 0x7630 */
            {8'h00}, /* 0x762f */
            {8'h00}, /* 0x762e */
            {8'h00}, /* 0x762d */
            {8'h00}, /* 0x762c */
            {8'h00}, /* 0x762b */
            {8'h00}, /* 0x762a */
            {8'h00}, /* 0x7629 */
            {8'h00}, /* 0x7628 */
            {8'h00}, /* 0x7627 */
            {8'h00}, /* 0x7626 */
            {8'h00}, /* 0x7625 */
            {8'h00}, /* 0x7624 */
            {8'h00}, /* 0x7623 */
            {8'h00}, /* 0x7622 */
            {8'h00}, /* 0x7621 */
            {8'h00}, /* 0x7620 */
            {8'h00}, /* 0x761f */
            {8'h00}, /* 0x761e */
            {8'h00}, /* 0x761d */
            {8'h00}, /* 0x761c */
            {8'h00}, /* 0x761b */
            {8'h00}, /* 0x761a */
            {8'h00}, /* 0x7619 */
            {8'h00}, /* 0x7618 */
            {8'h00}, /* 0x7617 */
            {8'h00}, /* 0x7616 */
            {8'h00}, /* 0x7615 */
            {8'h00}, /* 0x7614 */
            {8'h00}, /* 0x7613 */
            {8'h00}, /* 0x7612 */
            {8'h00}, /* 0x7611 */
            {8'h00}, /* 0x7610 */
            {8'h00}, /* 0x760f */
            {8'h00}, /* 0x760e */
            {8'h00}, /* 0x760d */
            {8'h00}, /* 0x760c */
            {8'h00}, /* 0x760b */
            {8'h00}, /* 0x760a */
            {8'h00}, /* 0x7609 */
            {8'h00}, /* 0x7608 */
            {8'h00}, /* 0x7607 */
            {8'h00}, /* 0x7606 */
            {8'h00}, /* 0x7605 */
            {8'h00}, /* 0x7604 */
            {8'h00}, /* 0x7603 */
            {8'h00}, /* 0x7602 */
            {8'h00}, /* 0x7601 */
            {8'h00}, /* 0x7600 */
            {8'h00}, /* 0x75ff */
            {8'h00}, /* 0x75fe */
            {8'h00}, /* 0x75fd */
            {8'h00}, /* 0x75fc */
            {8'h00}, /* 0x75fb */
            {8'h00}, /* 0x75fa */
            {8'h00}, /* 0x75f9 */
            {8'h00}, /* 0x75f8 */
            {8'h00}, /* 0x75f7 */
            {8'h00}, /* 0x75f6 */
            {8'h00}, /* 0x75f5 */
            {8'h00}, /* 0x75f4 */
            {8'h00}, /* 0x75f3 */
            {8'h00}, /* 0x75f2 */
            {8'h00}, /* 0x75f1 */
            {8'h00}, /* 0x75f0 */
            {8'h00}, /* 0x75ef */
            {8'h00}, /* 0x75ee */
            {8'h00}, /* 0x75ed */
            {8'h00}, /* 0x75ec */
            {8'h00}, /* 0x75eb */
            {8'h00}, /* 0x75ea */
            {8'h00}, /* 0x75e9 */
            {8'h00}, /* 0x75e8 */
            {8'h00}, /* 0x75e7 */
            {8'h00}, /* 0x75e6 */
            {8'h00}, /* 0x75e5 */
            {8'h00}, /* 0x75e4 */
            {8'h00}, /* 0x75e3 */
            {8'h00}, /* 0x75e2 */
            {8'h00}, /* 0x75e1 */
            {8'h00}, /* 0x75e0 */
            {8'h00}, /* 0x75df */
            {8'h00}, /* 0x75de */
            {8'h00}, /* 0x75dd */
            {8'h00}, /* 0x75dc */
            {8'h00}, /* 0x75db */
            {8'h00}, /* 0x75da */
            {8'h00}, /* 0x75d9 */
            {8'h00}, /* 0x75d8 */
            {8'h00}, /* 0x75d7 */
            {8'h00}, /* 0x75d6 */
            {8'h00}, /* 0x75d5 */
            {8'h00}, /* 0x75d4 */
            {8'h00}, /* 0x75d3 */
            {8'h00}, /* 0x75d2 */
            {8'h00}, /* 0x75d1 */
            {8'h00}, /* 0x75d0 */
            {8'h00}, /* 0x75cf */
            {8'h00}, /* 0x75ce */
            {8'h00}, /* 0x75cd */
            {8'h00}, /* 0x75cc */
            {8'h00}, /* 0x75cb */
            {8'h00}, /* 0x75ca */
            {8'h00}, /* 0x75c9 */
            {8'h00}, /* 0x75c8 */
            {8'h00}, /* 0x75c7 */
            {8'h00}, /* 0x75c6 */
            {8'h00}, /* 0x75c5 */
            {8'h00}, /* 0x75c4 */
            {8'h00}, /* 0x75c3 */
            {8'h00}, /* 0x75c2 */
            {8'h00}, /* 0x75c1 */
            {8'h00}, /* 0x75c0 */
            {8'h00}, /* 0x75bf */
            {8'h00}, /* 0x75be */
            {8'h00}, /* 0x75bd */
            {8'h00}, /* 0x75bc */
            {8'h00}, /* 0x75bb */
            {8'h00}, /* 0x75ba */
            {8'h00}, /* 0x75b9 */
            {8'h00}, /* 0x75b8 */
            {8'h00}, /* 0x75b7 */
            {8'h00}, /* 0x75b6 */
            {8'h00}, /* 0x75b5 */
            {8'h00}, /* 0x75b4 */
            {8'h00}, /* 0x75b3 */
            {8'h00}, /* 0x75b2 */
            {8'h00}, /* 0x75b1 */
            {8'h00}, /* 0x75b0 */
            {8'h00}, /* 0x75af */
            {8'h00}, /* 0x75ae */
            {8'h00}, /* 0x75ad */
            {8'h00}, /* 0x75ac */
            {8'h00}, /* 0x75ab */
            {8'h00}, /* 0x75aa */
            {8'h00}, /* 0x75a9 */
            {8'h00}, /* 0x75a8 */
            {8'h00}, /* 0x75a7 */
            {8'h00}, /* 0x75a6 */
            {8'h00}, /* 0x75a5 */
            {8'h00}, /* 0x75a4 */
            {8'h00}, /* 0x75a3 */
            {8'h00}, /* 0x75a2 */
            {8'h00}, /* 0x75a1 */
            {8'h00}, /* 0x75a0 */
            {8'h00}, /* 0x759f */
            {8'h00}, /* 0x759e */
            {8'h00}, /* 0x759d */
            {8'h00}, /* 0x759c */
            {8'h00}, /* 0x759b */
            {8'h00}, /* 0x759a */
            {8'h00}, /* 0x7599 */
            {8'h00}, /* 0x7598 */
            {8'h00}, /* 0x7597 */
            {8'h00}, /* 0x7596 */
            {8'h00}, /* 0x7595 */
            {8'h00}, /* 0x7594 */
            {8'h00}, /* 0x7593 */
            {8'h00}, /* 0x7592 */
            {8'h00}, /* 0x7591 */
            {8'h00}, /* 0x7590 */
            {8'h00}, /* 0x758f */
            {8'h00}, /* 0x758e */
            {8'h00}, /* 0x758d */
            {8'h00}, /* 0x758c */
            {8'h00}, /* 0x758b */
            {8'h00}, /* 0x758a */
            {8'h00}, /* 0x7589 */
            {8'h00}, /* 0x7588 */
            {8'h00}, /* 0x7587 */
            {8'h00}, /* 0x7586 */
            {8'h00}, /* 0x7585 */
            {8'h00}, /* 0x7584 */
            {8'h00}, /* 0x7583 */
            {8'h00}, /* 0x7582 */
            {8'h00}, /* 0x7581 */
            {8'h00}, /* 0x7580 */
            {8'h00}, /* 0x757f */
            {8'h00}, /* 0x757e */
            {8'h00}, /* 0x757d */
            {8'h00}, /* 0x757c */
            {8'h00}, /* 0x757b */
            {8'h00}, /* 0x757a */
            {8'h00}, /* 0x7579 */
            {8'h00}, /* 0x7578 */
            {8'h00}, /* 0x7577 */
            {8'h00}, /* 0x7576 */
            {8'h00}, /* 0x7575 */
            {8'h00}, /* 0x7574 */
            {8'h00}, /* 0x7573 */
            {8'h00}, /* 0x7572 */
            {8'h00}, /* 0x7571 */
            {8'h00}, /* 0x7570 */
            {8'h00}, /* 0x756f */
            {8'h00}, /* 0x756e */
            {8'h00}, /* 0x756d */
            {8'h00}, /* 0x756c */
            {8'h00}, /* 0x756b */
            {8'h00}, /* 0x756a */
            {8'h00}, /* 0x7569 */
            {8'h00}, /* 0x7568 */
            {8'h00}, /* 0x7567 */
            {8'h00}, /* 0x7566 */
            {8'h00}, /* 0x7565 */
            {8'h00}, /* 0x7564 */
            {8'h00}, /* 0x7563 */
            {8'h00}, /* 0x7562 */
            {8'h00}, /* 0x7561 */
            {8'h00}, /* 0x7560 */
            {8'h00}, /* 0x755f */
            {8'h00}, /* 0x755e */
            {8'h00}, /* 0x755d */
            {8'h00}, /* 0x755c */
            {8'h00}, /* 0x755b */
            {8'h00}, /* 0x755a */
            {8'h00}, /* 0x7559 */
            {8'h00}, /* 0x7558 */
            {8'h00}, /* 0x7557 */
            {8'h00}, /* 0x7556 */
            {8'h00}, /* 0x7555 */
            {8'h00}, /* 0x7554 */
            {8'h00}, /* 0x7553 */
            {8'h00}, /* 0x7552 */
            {8'h00}, /* 0x7551 */
            {8'h00}, /* 0x7550 */
            {8'h00}, /* 0x754f */
            {8'h00}, /* 0x754e */
            {8'h00}, /* 0x754d */
            {8'h00}, /* 0x754c */
            {8'h00}, /* 0x754b */
            {8'h00}, /* 0x754a */
            {8'h00}, /* 0x7549 */
            {8'h00}, /* 0x7548 */
            {8'h00}, /* 0x7547 */
            {8'h00}, /* 0x7546 */
            {8'h00}, /* 0x7545 */
            {8'h00}, /* 0x7544 */
            {8'h00}, /* 0x7543 */
            {8'h00}, /* 0x7542 */
            {8'h00}, /* 0x7541 */
            {8'h00}, /* 0x7540 */
            {8'h00}, /* 0x753f */
            {8'h00}, /* 0x753e */
            {8'h00}, /* 0x753d */
            {8'h00}, /* 0x753c */
            {8'h00}, /* 0x753b */
            {8'h00}, /* 0x753a */
            {8'h00}, /* 0x7539 */
            {8'h00}, /* 0x7538 */
            {8'h00}, /* 0x7537 */
            {8'h00}, /* 0x7536 */
            {8'h00}, /* 0x7535 */
            {8'h00}, /* 0x7534 */
            {8'h00}, /* 0x7533 */
            {8'h00}, /* 0x7532 */
            {8'h00}, /* 0x7531 */
            {8'h00}, /* 0x7530 */
            {8'h00}, /* 0x752f */
            {8'h00}, /* 0x752e */
            {8'h00}, /* 0x752d */
            {8'h00}, /* 0x752c */
            {8'h00}, /* 0x752b */
            {8'h00}, /* 0x752a */
            {8'h00}, /* 0x7529 */
            {8'h00}, /* 0x7528 */
            {8'h00}, /* 0x7527 */
            {8'h00}, /* 0x7526 */
            {8'h00}, /* 0x7525 */
            {8'h00}, /* 0x7524 */
            {8'h00}, /* 0x7523 */
            {8'h00}, /* 0x7522 */
            {8'h00}, /* 0x7521 */
            {8'h00}, /* 0x7520 */
            {8'h00}, /* 0x751f */
            {8'h00}, /* 0x751e */
            {8'h00}, /* 0x751d */
            {8'h00}, /* 0x751c */
            {8'h00}, /* 0x751b */
            {8'h00}, /* 0x751a */
            {8'h00}, /* 0x7519 */
            {8'h00}, /* 0x7518 */
            {8'h00}, /* 0x7517 */
            {8'h00}, /* 0x7516 */
            {8'h00}, /* 0x7515 */
            {8'h00}, /* 0x7514 */
            {8'h00}, /* 0x7513 */
            {8'h00}, /* 0x7512 */
            {8'h00}, /* 0x7511 */
            {8'h00}, /* 0x7510 */
            {8'h00}, /* 0x750f */
            {8'h00}, /* 0x750e */
            {8'h00}, /* 0x750d */
            {8'h00}, /* 0x750c */
            {8'h00}, /* 0x750b */
            {8'h00}, /* 0x750a */
            {8'h00}, /* 0x7509 */
            {8'h00}, /* 0x7508 */
            {8'h00}, /* 0x7507 */
            {8'h00}, /* 0x7506 */
            {8'h00}, /* 0x7505 */
            {8'h00}, /* 0x7504 */
            {8'h00}, /* 0x7503 */
            {8'h00}, /* 0x7502 */
            {8'h00}, /* 0x7501 */
            {8'h00}, /* 0x7500 */
            {8'h00}, /* 0x74ff */
            {8'h00}, /* 0x74fe */
            {8'h00}, /* 0x74fd */
            {8'h00}, /* 0x74fc */
            {8'h00}, /* 0x74fb */
            {8'h00}, /* 0x74fa */
            {8'h00}, /* 0x74f9 */
            {8'h00}, /* 0x74f8 */
            {8'h00}, /* 0x74f7 */
            {8'h00}, /* 0x74f6 */
            {8'h00}, /* 0x74f5 */
            {8'h00}, /* 0x74f4 */
            {8'h00}, /* 0x74f3 */
            {8'h00}, /* 0x74f2 */
            {8'h00}, /* 0x74f1 */
            {8'h00}, /* 0x74f0 */
            {8'h00}, /* 0x74ef */
            {8'h00}, /* 0x74ee */
            {8'h00}, /* 0x74ed */
            {8'h00}, /* 0x74ec */
            {8'h00}, /* 0x74eb */
            {8'h00}, /* 0x74ea */
            {8'h00}, /* 0x74e9 */
            {8'h00}, /* 0x74e8 */
            {8'h00}, /* 0x74e7 */
            {8'h00}, /* 0x74e6 */
            {8'h00}, /* 0x74e5 */
            {8'h00}, /* 0x74e4 */
            {8'h00}, /* 0x74e3 */
            {8'h00}, /* 0x74e2 */
            {8'h00}, /* 0x74e1 */
            {8'h00}, /* 0x74e0 */
            {8'h00}, /* 0x74df */
            {8'h00}, /* 0x74de */
            {8'h00}, /* 0x74dd */
            {8'h00}, /* 0x74dc */
            {8'h00}, /* 0x74db */
            {8'h00}, /* 0x74da */
            {8'h00}, /* 0x74d9 */
            {8'h00}, /* 0x74d8 */
            {8'h00}, /* 0x74d7 */
            {8'h00}, /* 0x74d6 */
            {8'h00}, /* 0x74d5 */
            {8'h00}, /* 0x74d4 */
            {8'h00}, /* 0x74d3 */
            {8'h00}, /* 0x74d2 */
            {8'h00}, /* 0x74d1 */
            {8'h00}, /* 0x74d0 */
            {8'h00}, /* 0x74cf */
            {8'h00}, /* 0x74ce */
            {8'h00}, /* 0x74cd */
            {8'h00}, /* 0x74cc */
            {8'h00}, /* 0x74cb */
            {8'h00}, /* 0x74ca */
            {8'h00}, /* 0x74c9 */
            {8'h00}, /* 0x74c8 */
            {8'h00}, /* 0x74c7 */
            {8'h00}, /* 0x74c6 */
            {8'h00}, /* 0x74c5 */
            {8'h00}, /* 0x74c4 */
            {8'h00}, /* 0x74c3 */
            {8'h00}, /* 0x74c2 */
            {8'h00}, /* 0x74c1 */
            {8'h00}, /* 0x74c0 */
            {8'h00}, /* 0x74bf */
            {8'h00}, /* 0x74be */
            {8'h00}, /* 0x74bd */
            {8'h00}, /* 0x74bc */
            {8'h00}, /* 0x74bb */
            {8'h00}, /* 0x74ba */
            {8'h00}, /* 0x74b9 */
            {8'h00}, /* 0x74b8 */
            {8'h00}, /* 0x74b7 */
            {8'h00}, /* 0x74b6 */
            {8'h00}, /* 0x74b5 */
            {8'h00}, /* 0x74b4 */
            {8'h00}, /* 0x74b3 */
            {8'h00}, /* 0x74b2 */
            {8'h00}, /* 0x74b1 */
            {8'h00}, /* 0x74b0 */
            {8'h00}, /* 0x74af */
            {8'h00}, /* 0x74ae */
            {8'h00}, /* 0x74ad */
            {8'h00}, /* 0x74ac */
            {8'h00}, /* 0x74ab */
            {8'h00}, /* 0x74aa */
            {8'h00}, /* 0x74a9 */
            {8'h00}, /* 0x74a8 */
            {8'h00}, /* 0x74a7 */
            {8'h00}, /* 0x74a6 */
            {8'h00}, /* 0x74a5 */
            {8'h00}, /* 0x74a4 */
            {8'h00}, /* 0x74a3 */
            {8'h00}, /* 0x74a2 */
            {8'h00}, /* 0x74a1 */
            {8'h00}, /* 0x74a0 */
            {8'h00}, /* 0x749f */
            {8'h00}, /* 0x749e */
            {8'h00}, /* 0x749d */
            {8'h00}, /* 0x749c */
            {8'h00}, /* 0x749b */
            {8'h00}, /* 0x749a */
            {8'h00}, /* 0x7499 */
            {8'h00}, /* 0x7498 */
            {8'h00}, /* 0x7497 */
            {8'h00}, /* 0x7496 */
            {8'h00}, /* 0x7495 */
            {8'h00}, /* 0x7494 */
            {8'h00}, /* 0x7493 */
            {8'h00}, /* 0x7492 */
            {8'h00}, /* 0x7491 */
            {8'h00}, /* 0x7490 */
            {8'h00}, /* 0x748f */
            {8'h00}, /* 0x748e */
            {8'h00}, /* 0x748d */
            {8'h00}, /* 0x748c */
            {8'h00}, /* 0x748b */
            {8'h00}, /* 0x748a */
            {8'h00}, /* 0x7489 */
            {8'h00}, /* 0x7488 */
            {8'h00}, /* 0x7487 */
            {8'h00}, /* 0x7486 */
            {8'h00}, /* 0x7485 */
            {8'h00}, /* 0x7484 */
            {8'h00}, /* 0x7483 */
            {8'h00}, /* 0x7482 */
            {8'h00}, /* 0x7481 */
            {8'h00}, /* 0x7480 */
            {8'h00}, /* 0x747f */
            {8'h00}, /* 0x747e */
            {8'h00}, /* 0x747d */
            {8'h00}, /* 0x747c */
            {8'h00}, /* 0x747b */
            {8'h00}, /* 0x747a */
            {8'h00}, /* 0x7479 */
            {8'h00}, /* 0x7478 */
            {8'h00}, /* 0x7477 */
            {8'h00}, /* 0x7476 */
            {8'h00}, /* 0x7475 */
            {8'h00}, /* 0x7474 */
            {8'h00}, /* 0x7473 */
            {8'h00}, /* 0x7472 */
            {8'h00}, /* 0x7471 */
            {8'h00}, /* 0x7470 */
            {8'h00}, /* 0x746f */
            {8'h00}, /* 0x746e */
            {8'h00}, /* 0x746d */
            {8'h00}, /* 0x746c */
            {8'h00}, /* 0x746b */
            {8'h00}, /* 0x746a */
            {8'h00}, /* 0x7469 */
            {8'h00}, /* 0x7468 */
            {8'h00}, /* 0x7467 */
            {8'h00}, /* 0x7466 */
            {8'h00}, /* 0x7465 */
            {8'h00}, /* 0x7464 */
            {8'h00}, /* 0x7463 */
            {8'h00}, /* 0x7462 */
            {8'h00}, /* 0x7461 */
            {8'h00}, /* 0x7460 */
            {8'h00}, /* 0x745f */
            {8'h00}, /* 0x745e */
            {8'h00}, /* 0x745d */
            {8'h00}, /* 0x745c */
            {8'h00}, /* 0x745b */
            {8'h00}, /* 0x745a */
            {8'h00}, /* 0x7459 */
            {8'h00}, /* 0x7458 */
            {8'h00}, /* 0x7457 */
            {8'h00}, /* 0x7456 */
            {8'h00}, /* 0x7455 */
            {8'h00}, /* 0x7454 */
            {8'h00}, /* 0x7453 */
            {8'h00}, /* 0x7452 */
            {8'h00}, /* 0x7451 */
            {8'h00}, /* 0x7450 */
            {8'h00}, /* 0x744f */
            {8'h00}, /* 0x744e */
            {8'h00}, /* 0x744d */
            {8'h00}, /* 0x744c */
            {8'h00}, /* 0x744b */
            {8'h00}, /* 0x744a */
            {8'h00}, /* 0x7449 */
            {8'h00}, /* 0x7448 */
            {8'h00}, /* 0x7447 */
            {8'h00}, /* 0x7446 */
            {8'h00}, /* 0x7445 */
            {8'h00}, /* 0x7444 */
            {8'h00}, /* 0x7443 */
            {8'h00}, /* 0x7442 */
            {8'h00}, /* 0x7441 */
            {8'h00}, /* 0x7440 */
            {8'h00}, /* 0x743f */
            {8'h00}, /* 0x743e */
            {8'h00}, /* 0x743d */
            {8'h00}, /* 0x743c */
            {8'h00}, /* 0x743b */
            {8'h00}, /* 0x743a */
            {8'h00}, /* 0x7439 */
            {8'h00}, /* 0x7438 */
            {8'h00}, /* 0x7437 */
            {8'h00}, /* 0x7436 */
            {8'h00}, /* 0x7435 */
            {8'h00}, /* 0x7434 */
            {8'h00}, /* 0x7433 */
            {8'h00}, /* 0x7432 */
            {8'h00}, /* 0x7431 */
            {8'h00}, /* 0x7430 */
            {8'h00}, /* 0x742f */
            {8'h00}, /* 0x742e */
            {8'h00}, /* 0x742d */
            {8'h00}, /* 0x742c */
            {8'h00}, /* 0x742b */
            {8'h00}, /* 0x742a */
            {8'h00}, /* 0x7429 */
            {8'h00}, /* 0x7428 */
            {8'h00}, /* 0x7427 */
            {8'h00}, /* 0x7426 */
            {8'h00}, /* 0x7425 */
            {8'h00}, /* 0x7424 */
            {8'h00}, /* 0x7423 */
            {8'h00}, /* 0x7422 */
            {8'h00}, /* 0x7421 */
            {8'h00}, /* 0x7420 */
            {8'h00}, /* 0x741f */
            {8'h00}, /* 0x741e */
            {8'h00}, /* 0x741d */
            {8'h00}, /* 0x741c */
            {8'h00}, /* 0x741b */
            {8'h00}, /* 0x741a */
            {8'h00}, /* 0x7419 */
            {8'h00}, /* 0x7418 */
            {8'h00}, /* 0x7417 */
            {8'h00}, /* 0x7416 */
            {8'h00}, /* 0x7415 */
            {8'h00}, /* 0x7414 */
            {8'h00}, /* 0x7413 */
            {8'h00}, /* 0x7412 */
            {8'h00}, /* 0x7411 */
            {8'h00}, /* 0x7410 */
            {8'h00}, /* 0x740f */
            {8'h00}, /* 0x740e */
            {8'h00}, /* 0x740d */
            {8'h00}, /* 0x740c */
            {8'h00}, /* 0x740b */
            {8'h00}, /* 0x740a */
            {8'h00}, /* 0x7409 */
            {8'h00}, /* 0x7408 */
            {8'h00}, /* 0x7407 */
            {8'h00}, /* 0x7406 */
            {8'h00}, /* 0x7405 */
            {8'h00}, /* 0x7404 */
            {8'h00}, /* 0x7403 */
            {8'h00}, /* 0x7402 */
            {8'h00}, /* 0x7401 */
            {8'h00}, /* 0x7400 */
            {8'h00}, /* 0x73ff */
            {8'h00}, /* 0x73fe */
            {8'h00}, /* 0x73fd */
            {8'h00}, /* 0x73fc */
            {8'h00}, /* 0x73fb */
            {8'h00}, /* 0x73fa */
            {8'h00}, /* 0x73f9 */
            {8'h00}, /* 0x73f8 */
            {8'h00}, /* 0x73f7 */
            {8'h00}, /* 0x73f6 */
            {8'h00}, /* 0x73f5 */
            {8'h00}, /* 0x73f4 */
            {8'h00}, /* 0x73f3 */
            {8'h00}, /* 0x73f2 */
            {8'h00}, /* 0x73f1 */
            {8'h00}, /* 0x73f0 */
            {8'h00}, /* 0x73ef */
            {8'h00}, /* 0x73ee */
            {8'h00}, /* 0x73ed */
            {8'h00}, /* 0x73ec */
            {8'h00}, /* 0x73eb */
            {8'h00}, /* 0x73ea */
            {8'h00}, /* 0x73e9 */
            {8'h00}, /* 0x73e8 */
            {8'h00}, /* 0x73e7 */
            {8'h00}, /* 0x73e6 */
            {8'h00}, /* 0x73e5 */
            {8'h00}, /* 0x73e4 */
            {8'h00}, /* 0x73e3 */
            {8'h00}, /* 0x73e2 */
            {8'h00}, /* 0x73e1 */
            {8'h00}, /* 0x73e0 */
            {8'h00}, /* 0x73df */
            {8'h00}, /* 0x73de */
            {8'h00}, /* 0x73dd */
            {8'h00}, /* 0x73dc */
            {8'h00}, /* 0x73db */
            {8'h00}, /* 0x73da */
            {8'h00}, /* 0x73d9 */
            {8'h00}, /* 0x73d8 */
            {8'h00}, /* 0x73d7 */
            {8'h00}, /* 0x73d6 */
            {8'h00}, /* 0x73d5 */
            {8'h00}, /* 0x73d4 */
            {8'h00}, /* 0x73d3 */
            {8'h00}, /* 0x73d2 */
            {8'h00}, /* 0x73d1 */
            {8'h00}, /* 0x73d0 */
            {8'h00}, /* 0x73cf */
            {8'h00}, /* 0x73ce */
            {8'h00}, /* 0x73cd */
            {8'h00}, /* 0x73cc */
            {8'h00}, /* 0x73cb */
            {8'h00}, /* 0x73ca */
            {8'h00}, /* 0x73c9 */
            {8'h00}, /* 0x73c8 */
            {8'h00}, /* 0x73c7 */
            {8'h00}, /* 0x73c6 */
            {8'h00}, /* 0x73c5 */
            {8'h00}, /* 0x73c4 */
            {8'h00}, /* 0x73c3 */
            {8'h00}, /* 0x73c2 */
            {8'h00}, /* 0x73c1 */
            {8'h00}, /* 0x73c0 */
            {8'h00}, /* 0x73bf */
            {8'h00}, /* 0x73be */
            {8'h00}, /* 0x73bd */
            {8'h00}, /* 0x73bc */
            {8'h00}, /* 0x73bb */
            {8'h00}, /* 0x73ba */
            {8'h00}, /* 0x73b9 */
            {8'h00}, /* 0x73b8 */
            {8'h00}, /* 0x73b7 */
            {8'h00}, /* 0x73b6 */
            {8'h00}, /* 0x73b5 */
            {8'h00}, /* 0x73b4 */
            {8'h00}, /* 0x73b3 */
            {8'h00}, /* 0x73b2 */
            {8'h00}, /* 0x73b1 */
            {8'h00}, /* 0x73b0 */
            {8'h00}, /* 0x73af */
            {8'h00}, /* 0x73ae */
            {8'h00}, /* 0x73ad */
            {8'h00}, /* 0x73ac */
            {8'h00}, /* 0x73ab */
            {8'h00}, /* 0x73aa */
            {8'h00}, /* 0x73a9 */
            {8'h00}, /* 0x73a8 */
            {8'h00}, /* 0x73a7 */
            {8'h00}, /* 0x73a6 */
            {8'h00}, /* 0x73a5 */
            {8'h00}, /* 0x73a4 */
            {8'h00}, /* 0x73a3 */
            {8'h00}, /* 0x73a2 */
            {8'h00}, /* 0x73a1 */
            {8'h00}, /* 0x73a0 */
            {8'h00}, /* 0x739f */
            {8'h00}, /* 0x739e */
            {8'h00}, /* 0x739d */
            {8'h00}, /* 0x739c */
            {8'h00}, /* 0x739b */
            {8'h00}, /* 0x739a */
            {8'h00}, /* 0x7399 */
            {8'h00}, /* 0x7398 */
            {8'h00}, /* 0x7397 */
            {8'h00}, /* 0x7396 */
            {8'h00}, /* 0x7395 */
            {8'h00}, /* 0x7394 */
            {8'h00}, /* 0x7393 */
            {8'h00}, /* 0x7392 */
            {8'h00}, /* 0x7391 */
            {8'h00}, /* 0x7390 */
            {8'h00}, /* 0x738f */
            {8'h00}, /* 0x738e */
            {8'h00}, /* 0x738d */
            {8'h00}, /* 0x738c */
            {8'h00}, /* 0x738b */
            {8'h00}, /* 0x738a */
            {8'h00}, /* 0x7389 */
            {8'h00}, /* 0x7388 */
            {8'h00}, /* 0x7387 */
            {8'h00}, /* 0x7386 */
            {8'h00}, /* 0x7385 */
            {8'h00}, /* 0x7384 */
            {8'h00}, /* 0x7383 */
            {8'h00}, /* 0x7382 */
            {8'h00}, /* 0x7381 */
            {8'h00}, /* 0x7380 */
            {8'h00}, /* 0x737f */
            {8'h00}, /* 0x737e */
            {8'h00}, /* 0x737d */
            {8'h00}, /* 0x737c */
            {8'h00}, /* 0x737b */
            {8'h00}, /* 0x737a */
            {8'h00}, /* 0x7379 */
            {8'h00}, /* 0x7378 */
            {8'h00}, /* 0x7377 */
            {8'h00}, /* 0x7376 */
            {8'h00}, /* 0x7375 */
            {8'h00}, /* 0x7374 */
            {8'h00}, /* 0x7373 */
            {8'h00}, /* 0x7372 */
            {8'h00}, /* 0x7371 */
            {8'h00}, /* 0x7370 */
            {8'h00}, /* 0x736f */
            {8'h00}, /* 0x736e */
            {8'h00}, /* 0x736d */
            {8'h00}, /* 0x736c */
            {8'h00}, /* 0x736b */
            {8'h00}, /* 0x736a */
            {8'h00}, /* 0x7369 */
            {8'h00}, /* 0x7368 */
            {8'h00}, /* 0x7367 */
            {8'h00}, /* 0x7366 */
            {8'h00}, /* 0x7365 */
            {8'h00}, /* 0x7364 */
            {8'h00}, /* 0x7363 */
            {8'h00}, /* 0x7362 */
            {8'h00}, /* 0x7361 */
            {8'h00}, /* 0x7360 */
            {8'h00}, /* 0x735f */
            {8'h00}, /* 0x735e */
            {8'h00}, /* 0x735d */
            {8'h00}, /* 0x735c */
            {8'h00}, /* 0x735b */
            {8'h00}, /* 0x735a */
            {8'h00}, /* 0x7359 */
            {8'h00}, /* 0x7358 */
            {8'h00}, /* 0x7357 */
            {8'h00}, /* 0x7356 */
            {8'h00}, /* 0x7355 */
            {8'h00}, /* 0x7354 */
            {8'h00}, /* 0x7353 */
            {8'h00}, /* 0x7352 */
            {8'h00}, /* 0x7351 */
            {8'h00}, /* 0x7350 */
            {8'h00}, /* 0x734f */
            {8'h00}, /* 0x734e */
            {8'h00}, /* 0x734d */
            {8'h00}, /* 0x734c */
            {8'h00}, /* 0x734b */
            {8'h00}, /* 0x734a */
            {8'h00}, /* 0x7349 */
            {8'h00}, /* 0x7348 */
            {8'h00}, /* 0x7347 */
            {8'h00}, /* 0x7346 */
            {8'h00}, /* 0x7345 */
            {8'h00}, /* 0x7344 */
            {8'h00}, /* 0x7343 */
            {8'h00}, /* 0x7342 */
            {8'h00}, /* 0x7341 */
            {8'h00}, /* 0x7340 */
            {8'h00}, /* 0x733f */
            {8'h00}, /* 0x733e */
            {8'h00}, /* 0x733d */
            {8'h00}, /* 0x733c */
            {8'h00}, /* 0x733b */
            {8'h00}, /* 0x733a */
            {8'h00}, /* 0x7339 */
            {8'h00}, /* 0x7338 */
            {8'h00}, /* 0x7337 */
            {8'h00}, /* 0x7336 */
            {8'h00}, /* 0x7335 */
            {8'h00}, /* 0x7334 */
            {8'h00}, /* 0x7333 */
            {8'h00}, /* 0x7332 */
            {8'h00}, /* 0x7331 */
            {8'h00}, /* 0x7330 */
            {8'h00}, /* 0x732f */
            {8'h00}, /* 0x732e */
            {8'h00}, /* 0x732d */
            {8'h00}, /* 0x732c */
            {8'h00}, /* 0x732b */
            {8'h00}, /* 0x732a */
            {8'h00}, /* 0x7329 */
            {8'h00}, /* 0x7328 */
            {8'h00}, /* 0x7327 */
            {8'h00}, /* 0x7326 */
            {8'h00}, /* 0x7325 */
            {8'h00}, /* 0x7324 */
            {8'h00}, /* 0x7323 */
            {8'h00}, /* 0x7322 */
            {8'h00}, /* 0x7321 */
            {8'h00}, /* 0x7320 */
            {8'h00}, /* 0x731f */
            {8'h00}, /* 0x731e */
            {8'h00}, /* 0x731d */
            {8'h00}, /* 0x731c */
            {8'h00}, /* 0x731b */
            {8'h00}, /* 0x731a */
            {8'h00}, /* 0x7319 */
            {8'h00}, /* 0x7318 */
            {8'h00}, /* 0x7317 */
            {8'h00}, /* 0x7316 */
            {8'h00}, /* 0x7315 */
            {8'h00}, /* 0x7314 */
            {8'h00}, /* 0x7313 */
            {8'h00}, /* 0x7312 */
            {8'h00}, /* 0x7311 */
            {8'h00}, /* 0x7310 */
            {8'h00}, /* 0x730f */
            {8'h00}, /* 0x730e */
            {8'h00}, /* 0x730d */
            {8'h00}, /* 0x730c */
            {8'h00}, /* 0x730b */
            {8'h00}, /* 0x730a */
            {8'h00}, /* 0x7309 */
            {8'h00}, /* 0x7308 */
            {8'h00}, /* 0x7307 */
            {8'h00}, /* 0x7306 */
            {8'h00}, /* 0x7305 */
            {8'h00}, /* 0x7304 */
            {8'h00}, /* 0x7303 */
            {8'h00}, /* 0x7302 */
            {8'h00}, /* 0x7301 */
            {8'h00}, /* 0x7300 */
            {8'h00}, /* 0x72ff */
            {8'h00}, /* 0x72fe */
            {8'h00}, /* 0x72fd */
            {8'h00}, /* 0x72fc */
            {8'h00}, /* 0x72fb */
            {8'h00}, /* 0x72fa */
            {8'h00}, /* 0x72f9 */
            {8'h00}, /* 0x72f8 */
            {8'h00}, /* 0x72f7 */
            {8'h00}, /* 0x72f6 */
            {8'h00}, /* 0x72f5 */
            {8'h00}, /* 0x72f4 */
            {8'h00}, /* 0x72f3 */
            {8'h00}, /* 0x72f2 */
            {8'h00}, /* 0x72f1 */
            {8'h00}, /* 0x72f0 */
            {8'h00}, /* 0x72ef */
            {8'h00}, /* 0x72ee */
            {8'h00}, /* 0x72ed */
            {8'h00}, /* 0x72ec */
            {8'h00}, /* 0x72eb */
            {8'h00}, /* 0x72ea */
            {8'h00}, /* 0x72e9 */
            {8'h00}, /* 0x72e8 */
            {8'h00}, /* 0x72e7 */
            {8'h00}, /* 0x72e6 */
            {8'h00}, /* 0x72e5 */
            {8'h00}, /* 0x72e4 */
            {8'h00}, /* 0x72e3 */
            {8'h00}, /* 0x72e2 */
            {8'h00}, /* 0x72e1 */
            {8'h00}, /* 0x72e0 */
            {8'h00}, /* 0x72df */
            {8'h00}, /* 0x72de */
            {8'h00}, /* 0x72dd */
            {8'h00}, /* 0x72dc */
            {8'h00}, /* 0x72db */
            {8'h00}, /* 0x72da */
            {8'h00}, /* 0x72d9 */
            {8'h00}, /* 0x72d8 */
            {8'h00}, /* 0x72d7 */
            {8'h00}, /* 0x72d6 */
            {8'h00}, /* 0x72d5 */
            {8'h00}, /* 0x72d4 */
            {8'h00}, /* 0x72d3 */
            {8'h00}, /* 0x72d2 */
            {8'h00}, /* 0x72d1 */
            {8'h00}, /* 0x72d0 */
            {8'h00}, /* 0x72cf */
            {8'h00}, /* 0x72ce */
            {8'h00}, /* 0x72cd */
            {8'h00}, /* 0x72cc */
            {8'h00}, /* 0x72cb */
            {8'h00}, /* 0x72ca */
            {8'h00}, /* 0x72c9 */
            {8'h00}, /* 0x72c8 */
            {8'h00}, /* 0x72c7 */
            {8'h00}, /* 0x72c6 */
            {8'h00}, /* 0x72c5 */
            {8'h00}, /* 0x72c4 */
            {8'h00}, /* 0x72c3 */
            {8'h00}, /* 0x72c2 */
            {8'h00}, /* 0x72c1 */
            {8'h00}, /* 0x72c0 */
            {8'h00}, /* 0x72bf */
            {8'h00}, /* 0x72be */
            {8'h00}, /* 0x72bd */
            {8'h00}, /* 0x72bc */
            {8'h00}, /* 0x72bb */
            {8'h00}, /* 0x72ba */
            {8'h00}, /* 0x72b9 */
            {8'h00}, /* 0x72b8 */
            {8'h00}, /* 0x72b7 */
            {8'h00}, /* 0x72b6 */
            {8'h00}, /* 0x72b5 */
            {8'h00}, /* 0x72b4 */
            {8'h00}, /* 0x72b3 */
            {8'h00}, /* 0x72b2 */
            {8'h00}, /* 0x72b1 */
            {8'h00}, /* 0x72b0 */
            {8'h00}, /* 0x72af */
            {8'h00}, /* 0x72ae */
            {8'h00}, /* 0x72ad */
            {8'h00}, /* 0x72ac */
            {8'h00}, /* 0x72ab */
            {8'h00}, /* 0x72aa */
            {8'h00}, /* 0x72a9 */
            {8'h00}, /* 0x72a8 */
            {8'h00}, /* 0x72a7 */
            {8'h00}, /* 0x72a6 */
            {8'h00}, /* 0x72a5 */
            {8'h00}, /* 0x72a4 */
            {8'h00}, /* 0x72a3 */
            {8'h00}, /* 0x72a2 */
            {8'h00}, /* 0x72a1 */
            {8'h00}, /* 0x72a0 */
            {8'h00}, /* 0x729f */
            {8'h00}, /* 0x729e */
            {8'h00}, /* 0x729d */
            {8'h00}, /* 0x729c */
            {8'h00}, /* 0x729b */
            {8'h00}, /* 0x729a */
            {8'h00}, /* 0x7299 */
            {8'h00}, /* 0x7298 */
            {8'h00}, /* 0x7297 */
            {8'h00}, /* 0x7296 */
            {8'h00}, /* 0x7295 */
            {8'h00}, /* 0x7294 */
            {8'h00}, /* 0x7293 */
            {8'h00}, /* 0x7292 */
            {8'h00}, /* 0x7291 */
            {8'h00}, /* 0x7290 */
            {8'h00}, /* 0x728f */
            {8'h00}, /* 0x728e */
            {8'h00}, /* 0x728d */
            {8'h00}, /* 0x728c */
            {8'h00}, /* 0x728b */
            {8'h00}, /* 0x728a */
            {8'h00}, /* 0x7289 */
            {8'h00}, /* 0x7288 */
            {8'h00}, /* 0x7287 */
            {8'h00}, /* 0x7286 */
            {8'h00}, /* 0x7285 */
            {8'h00}, /* 0x7284 */
            {8'h00}, /* 0x7283 */
            {8'h00}, /* 0x7282 */
            {8'h00}, /* 0x7281 */
            {8'h00}, /* 0x7280 */
            {8'h00}, /* 0x727f */
            {8'h00}, /* 0x727e */
            {8'h00}, /* 0x727d */
            {8'h00}, /* 0x727c */
            {8'h00}, /* 0x727b */
            {8'h00}, /* 0x727a */
            {8'h00}, /* 0x7279 */
            {8'h00}, /* 0x7278 */
            {8'h00}, /* 0x7277 */
            {8'h00}, /* 0x7276 */
            {8'h00}, /* 0x7275 */
            {8'h00}, /* 0x7274 */
            {8'h00}, /* 0x7273 */
            {8'h00}, /* 0x7272 */
            {8'h00}, /* 0x7271 */
            {8'h00}, /* 0x7270 */
            {8'h00}, /* 0x726f */
            {8'h00}, /* 0x726e */
            {8'h00}, /* 0x726d */
            {8'h00}, /* 0x726c */
            {8'h00}, /* 0x726b */
            {8'h00}, /* 0x726a */
            {8'h00}, /* 0x7269 */
            {8'h00}, /* 0x7268 */
            {8'h00}, /* 0x7267 */
            {8'h00}, /* 0x7266 */
            {8'h00}, /* 0x7265 */
            {8'h00}, /* 0x7264 */
            {8'h00}, /* 0x7263 */
            {8'h00}, /* 0x7262 */
            {8'h00}, /* 0x7261 */
            {8'h00}, /* 0x7260 */
            {8'h00}, /* 0x725f */
            {8'h00}, /* 0x725e */
            {8'h00}, /* 0x725d */
            {8'h00}, /* 0x725c */
            {8'h00}, /* 0x725b */
            {8'h00}, /* 0x725a */
            {8'h00}, /* 0x7259 */
            {8'h00}, /* 0x7258 */
            {8'h00}, /* 0x7257 */
            {8'h00}, /* 0x7256 */
            {8'h00}, /* 0x7255 */
            {8'h00}, /* 0x7254 */
            {8'h00}, /* 0x7253 */
            {8'h00}, /* 0x7252 */
            {8'h00}, /* 0x7251 */
            {8'h00}, /* 0x7250 */
            {8'h00}, /* 0x724f */
            {8'h00}, /* 0x724e */
            {8'h00}, /* 0x724d */
            {8'h00}, /* 0x724c */
            {8'h00}, /* 0x724b */
            {8'h00}, /* 0x724a */
            {8'h00}, /* 0x7249 */
            {8'h00}, /* 0x7248 */
            {8'h00}, /* 0x7247 */
            {8'h00}, /* 0x7246 */
            {8'h00}, /* 0x7245 */
            {8'h00}, /* 0x7244 */
            {8'h00}, /* 0x7243 */
            {8'h00}, /* 0x7242 */
            {8'h00}, /* 0x7241 */
            {8'h00}, /* 0x7240 */
            {8'h00}, /* 0x723f */
            {8'h00}, /* 0x723e */
            {8'h00}, /* 0x723d */
            {8'h00}, /* 0x723c */
            {8'h00}, /* 0x723b */
            {8'h00}, /* 0x723a */
            {8'h00}, /* 0x7239 */
            {8'h00}, /* 0x7238 */
            {8'h00}, /* 0x7237 */
            {8'h00}, /* 0x7236 */
            {8'h00}, /* 0x7235 */
            {8'h00}, /* 0x7234 */
            {8'h00}, /* 0x7233 */
            {8'h00}, /* 0x7232 */
            {8'h00}, /* 0x7231 */
            {8'h00}, /* 0x7230 */
            {8'h00}, /* 0x722f */
            {8'h00}, /* 0x722e */
            {8'h00}, /* 0x722d */
            {8'h00}, /* 0x722c */
            {8'h00}, /* 0x722b */
            {8'h00}, /* 0x722a */
            {8'h00}, /* 0x7229 */
            {8'h00}, /* 0x7228 */
            {8'h00}, /* 0x7227 */
            {8'h00}, /* 0x7226 */
            {8'h00}, /* 0x7225 */
            {8'h00}, /* 0x7224 */
            {8'h00}, /* 0x7223 */
            {8'h00}, /* 0x7222 */
            {8'h00}, /* 0x7221 */
            {8'h00}, /* 0x7220 */
            {8'h00}, /* 0x721f */
            {8'h00}, /* 0x721e */
            {8'h00}, /* 0x721d */
            {8'h00}, /* 0x721c */
            {8'h00}, /* 0x721b */
            {8'h00}, /* 0x721a */
            {8'h00}, /* 0x7219 */
            {8'h00}, /* 0x7218 */
            {8'h00}, /* 0x7217 */
            {8'h00}, /* 0x7216 */
            {8'h00}, /* 0x7215 */
            {8'h00}, /* 0x7214 */
            {8'h00}, /* 0x7213 */
            {8'h00}, /* 0x7212 */
            {8'h00}, /* 0x7211 */
            {8'h00}, /* 0x7210 */
            {8'h00}, /* 0x720f */
            {8'h00}, /* 0x720e */
            {8'h00}, /* 0x720d */
            {8'h00}, /* 0x720c */
            {8'h00}, /* 0x720b */
            {8'h00}, /* 0x720a */
            {8'h00}, /* 0x7209 */
            {8'h00}, /* 0x7208 */
            {8'h00}, /* 0x7207 */
            {8'h00}, /* 0x7206 */
            {8'h00}, /* 0x7205 */
            {8'h00}, /* 0x7204 */
            {8'h00}, /* 0x7203 */
            {8'h00}, /* 0x7202 */
            {8'h00}, /* 0x7201 */
            {8'h00}, /* 0x7200 */
            {8'h00}, /* 0x71ff */
            {8'h00}, /* 0x71fe */
            {8'h00}, /* 0x71fd */
            {8'h00}, /* 0x71fc */
            {8'h00}, /* 0x71fb */
            {8'h00}, /* 0x71fa */
            {8'h00}, /* 0x71f9 */
            {8'h00}, /* 0x71f8 */
            {8'h00}, /* 0x71f7 */
            {8'h00}, /* 0x71f6 */
            {8'h00}, /* 0x71f5 */
            {8'h00}, /* 0x71f4 */
            {8'h00}, /* 0x71f3 */
            {8'h00}, /* 0x71f2 */
            {8'h00}, /* 0x71f1 */
            {8'h00}, /* 0x71f0 */
            {8'h00}, /* 0x71ef */
            {8'h00}, /* 0x71ee */
            {8'h00}, /* 0x71ed */
            {8'h00}, /* 0x71ec */
            {8'h00}, /* 0x71eb */
            {8'h00}, /* 0x71ea */
            {8'h00}, /* 0x71e9 */
            {8'h00}, /* 0x71e8 */
            {8'h00}, /* 0x71e7 */
            {8'h00}, /* 0x71e6 */
            {8'h00}, /* 0x71e5 */
            {8'h00}, /* 0x71e4 */
            {8'h00}, /* 0x71e3 */
            {8'h00}, /* 0x71e2 */
            {8'h00}, /* 0x71e1 */
            {8'h00}, /* 0x71e0 */
            {8'h00}, /* 0x71df */
            {8'h00}, /* 0x71de */
            {8'h00}, /* 0x71dd */
            {8'h00}, /* 0x71dc */
            {8'h00}, /* 0x71db */
            {8'h00}, /* 0x71da */
            {8'h00}, /* 0x71d9 */
            {8'h00}, /* 0x71d8 */
            {8'h00}, /* 0x71d7 */
            {8'h00}, /* 0x71d6 */
            {8'h00}, /* 0x71d5 */
            {8'h00}, /* 0x71d4 */
            {8'h00}, /* 0x71d3 */
            {8'h00}, /* 0x71d2 */
            {8'h00}, /* 0x71d1 */
            {8'h00}, /* 0x71d0 */
            {8'h00}, /* 0x71cf */
            {8'h00}, /* 0x71ce */
            {8'h00}, /* 0x71cd */
            {8'h00}, /* 0x71cc */
            {8'h00}, /* 0x71cb */
            {8'h00}, /* 0x71ca */
            {8'h00}, /* 0x71c9 */
            {8'h00}, /* 0x71c8 */
            {8'h00}, /* 0x71c7 */
            {8'h00}, /* 0x71c6 */
            {8'h00}, /* 0x71c5 */
            {8'h00}, /* 0x71c4 */
            {8'h00}, /* 0x71c3 */
            {8'h00}, /* 0x71c2 */
            {8'h00}, /* 0x71c1 */
            {8'h00}, /* 0x71c0 */
            {8'h00}, /* 0x71bf */
            {8'h00}, /* 0x71be */
            {8'h00}, /* 0x71bd */
            {8'h00}, /* 0x71bc */
            {8'h00}, /* 0x71bb */
            {8'h00}, /* 0x71ba */
            {8'h00}, /* 0x71b9 */
            {8'h00}, /* 0x71b8 */
            {8'h00}, /* 0x71b7 */
            {8'h00}, /* 0x71b6 */
            {8'h00}, /* 0x71b5 */
            {8'h00}, /* 0x71b4 */
            {8'h00}, /* 0x71b3 */
            {8'h00}, /* 0x71b2 */
            {8'h00}, /* 0x71b1 */
            {8'h00}, /* 0x71b0 */
            {8'h00}, /* 0x71af */
            {8'h00}, /* 0x71ae */
            {8'h00}, /* 0x71ad */
            {8'h00}, /* 0x71ac */
            {8'h00}, /* 0x71ab */
            {8'h00}, /* 0x71aa */
            {8'h00}, /* 0x71a9 */
            {8'h00}, /* 0x71a8 */
            {8'h00}, /* 0x71a7 */
            {8'h00}, /* 0x71a6 */
            {8'h00}, /* 0x71a5 */
            {8'h00}, /* 0x71a4 */
            {8'h00}, /* 0x71a3 */
            {8'h00}, /* 0x71a2 */
            {8'h00}, /* 0x71a1 */
            {8'h00}, /* 0x71a0 */
            {8'h00}, /* 0x719f */
            {8'h00}, /* 0x719e */
            {8'h00}, /* 0x719d */
            {8'h00}, /* 0x719c */
            {8'h00}, /* 0x719b */
            {8'h00}, /* 0x719a */
            {8'h00}, /* 0x7199 */
            {8'h00}, /* 0x7198 */
            {8'h00}, /* 0x7197 */
            {8'h00}, /* 0x7196 */
            {8'h00}, /* 0x7195 */
            {8'h00}, /* 0x7194 */
            {8'h00}, /* 0x7193 */
            {8'h00}, /* 0x7192 */
            {8'h00}, /* 0x7191 */
            {8'h00}, /* 0x7190 */
            {8'h00}, /* 0x718f */
            {8'h00}, /* 0x718e */
            {8'h00}, /* 0x718d */
            {8'h00}, /* 0x718c */
            {8'h00}, /* 0x718b */
            {8'h00}, /* 0x718a */
            {8'h00}, /* 0x7189 */
            {8'h00}, /* 0x7188 */
            {8'h00}, /* 0x7187 */
            {8'h00}, /* 0x7186 */
            {8'h00}, /* 0x7185 */
            {8'h00}, /* 0x7184 */
            {8'h00}, /* 0x7183 */
            {8'h00}, /* 0x7182 */
            {8'h00}, /* 0x7181 */
            {8'h00}, /* 0x7180 */
            {8'h00}, /* 0x717f */
            {8'h00}, /* 0x717e */
            {8'h00}, /* 0x717d */
            {8'h00}, /* 0x717c */
            {8'h00}, /* 0x717b */
            {8'h00}, /* 0x717a */
            {8'h00}, /* 0x7179 */
            {8'h00}, /* 0x7178 */
            {8'h00}, /* 0x7177 */
            {8'h00}, /* 0x7176 */
            {8'h00}, /* 0x7175 */
            {8'h00}, /* 0x7174 */
            {8'h00}, /* 0x7173 */
            {8'h00}, /* 0x7172 */
            {8'h00}, /* 0x7171 */
            {8'h00}, /* 0x7170 */
            {8'h00}, /* 0x716f */
            {8'h00}, /* 0x716e */
            {8'h00}, /* 0x716d */
            {8'h00}, /* 0x716c */
            {8'h00}, /* 0x716b */
            {8'h00}, /* 0x716a */
            {8'h00}, /* 0x7169 */
            {8'h00}, /* 0x7168 */
            {8'h00}, /* 0x7167 */
            {8'h00}, /* 0x7166 */
            {8'h00}, /* 0x7165 */
            {8'h00}, /* 0x7164 */
            {8'h00}, /* 0x7163 */
            {8'h00}, /* 0x7162 */
            {8'h00}, /* 0x7161 */
            {8'h00}, /* 0x7160 */
            {8'h00}, /* 0x715f */
            {8'h00}, /* 0x715e */
            {8'h00}, /* 0x715d */
            {8'h00}, /* 0x715c */
            {8'h00}, /* 0x715b */
            {8'h00}, /* 0x715a */
            {8'h00}, /* 0x7159 */
            {8'h00}, /* 0x7158 */
            {8'h00}, /* 0x7157 */
            {8'h00}, /* 0x7156 */
            {8'h00}, /* 0x7155 */
            {8'h00}, /* 0x7154 */
            {8'h00}, /* 0x7153 */
            {8'h00}, /* 0x7152 */
            {8'h00}, /* 0x7151 */
            {8'h00}, /* 0x7150 */
            {8'h00}, /* 0x714f */
            {8'h00}, /* 0x714e */
            {8'h00}, /* 0x714d */
            {8'h00}, /* 0x714c */
            {8'h00}, /* 0x714b */
            {8'h00}, /* 0x714a */
            {8'h00}, /* 0x7149 */
            {8'h00}, /* 0x7148 */
            {8'h00}, /* 0x7147 */
            {8'h00}, /* 0x7146 */
            {8'h00}, /* 0x7145 */
            {8'h00}, /* 0x7144 */
            {8'h00}, /* 0x7143 */
            {8'h00}, /* 0x7142 */
            {8'h00}, /* 0x7141 */
            {8'h00}, /* 0x7140 */
            {8'h00}, /* 0x713f */
            {8'h00}, /* 0x713e */
            {8'h00}, /* 0x713d */
            {8'h00}, /* 0x713c */
            {8'h00}, /* 0x713b */
            {8'h00}, /* 0x713a */
            {8'h00}, /* 0x7139 */
            {8'h00}, /* 0x7138 */
            {8'h00}, /* 0x7137 */
            {8'h00}, /* 0x7136 */
            {8'h00}, /* 0x7135 */
            {8'h00}, /* 0x7134 */
            {8'h00}, /* 0x7133 */
            {8'h00}, /* 0x7132 */
            {8'h00}, /* 0x7131 */
            {8'h00}, /* 0x7130 */
            {8'h00}, /* 0x712f */
            {8'h00}, /* 0x712e */
            {8'h00}, /* 0x712d */
            {8'h00}, /* 0x712c */
            {8'h00}, /* 0x712b */
            {8'h00}, /* 0x712a */
            {8'h00}, /* 0x7129 */
            {8'h00}, /* 0x7128 */
            {8'h00}, /* 0x7127 */
            {8'h00}, /* 0x7126 */
            {8'h00}, /* 0x7125 */
            {8'h00}, /* 0x7124 */
            {8'h00}, /* 0x7123 */
            {8'h00}, /* 0x7122 */
            {8'h00}, /* 0x7121 */
            {8'h00}, /* 0x7120 */
            {8'h00}, /* 0x711f */
            {8'h00}, /* 0x711e */
            {8'h00}, /* 0x711d */
            {8'h00}, /* 0x711c */
            {8'h00}, /* 0x711b */
            {8'h00}, /* 0x711a */
            {8'h00}, /* 0x7119 */
            {8'h00}, /* 0x7118 */
            {8'h00}, /* 0x7117 */
            {8'h00}, /* 0x7116 */
            {8'h00}, /* 0x7115 */
            {8'h00}, /* 0x7114 */
            {8'h00}, /* 0x7113 */
            {8'h00}, /* 0x7112 */
            {8'h00}, /* 0x7111 */
            {8'h00}, /* 0x7110 */
            {8'h00}, /* 0x710f */
            {8'h00}, /* 0x710e */
            {8'h00}, /* 0x710d */
            {8'h00}, /* 0x710c */
            {8'h00}, /* 0x710b */
            {8'h00}, /* 0x710a */
            {8'h00}, /* 0x7109 */
            {8'h00}, /* 0x7108 */
            {8'h00}, /* 0x7107 */
            {8'h00}, /* 0x7106 */
            {8'h00}, /* 0x7105 */
            {8'h00}, /* 0x7104 */
            {8'h00}, /* 0x7103 */
            {8'h00}, /* 0x7102 */
            {8'h00}, /* 0x7101 */
            {8'h00}, /* 0x7100 */
            {8'h00}, /* 0x70ff */
            {8'h00}, /* 0x70fe */
            {8'h00}, /* 0x70fd */
            {8'h00}, /* 0x70fc */
            {8'h00}, /* 0x70fb */
            {8'h00}, /* 0x70fa */
            {8'h00}, /* 0x70f9 */
            {8'h00}, /* 0x70f8 */
            {8'h00}, /* 0x70f7 */
            {8'h00}, /* 0x70f6 */
            {8'h00}, /* 0x70f5 */
            {8'h00}, /* 0x70f4 */
            {8'h00}, /* 0x70f3 */
            {8'h00}, /* 0x70f2 */
            {8'h00}, /* 0x70f1 */
            {8'h00}, /* 0x70f0 */
            {8'h00}, /* 0x70ef */
            {8'h00}, /* 0x70ee */
            {8'h00}, /* 0x70ed */
            {8'h00}, /* 0x70ec */
            {8'h00}, /* 0x70eb */
            {8'h00}, /* 0x70ea */
            {8'h00}, /* 0x70e9 */
            {8'h00}, /* 0x70e8 */
            {8'h00}, /* 0x70e7 */
            {8'h00}, /* 0x70e6 */
            {8'h00}, /* 0x70e5 */
            {8'h00}, /* 0x70e4 */
            {8'h00}, /* 0x70e3 */
            {8'h00}, /* 0x70e2 */
            {8'h00}, /* 0x70e1 */
            {8'h00}, /* 0x70e0 */
            {8'h00}, /* 0x70df */
            {8'h00}, /* 0x70de */
            {8'h00}, /* 0x70dd */
            {8'h00}, /* 0x70dc */
            {8'h00}, /* 0x70db */
            {8'h00}, /* 0x70da */
            {8'h00}, /* 0x70d9 */
            {8'h00}, /* 0x70d8 */
            {8'h00}, /* 0x70d7 */
            {8'h00}, /* 0x70d6 */
            {8'h00}, /* 0x70d5 */
            {8'h00}, /* 0x70d4 */
            {8'h00}, /* 0x70d3 */
            {8'h00}, /* 0x70d2 */
            {8'h00}, /* 0x70d1 */
            {8'h00}, /* 0x70d0 */
            {8'h00}, /* 0x70cf */
            {8'h00}, /* 0x70ce */
            {8'h00}, /* 0x70cd */
            {8'h00}, /* 0x70cc */
            {8'h00}, /* 0x70cb */
            {8'h00}, /* 0x70ca */
            {8'h00}, /* 0x70c9 */
            {8'h00}, /* 0x70c8 */
            {8'h00}, /* 0x70c7 */
            {8'h00}, /* 0x70c6 */
            {8'h00}, /* 0x70c5 */
            {8'h00}, /* 0x70c4 */
            {8'h00}, /* 0x70c3 */
            {8'h00}, /* 0x70c2 */
            {8'h00}, /* 0x70c1 */
            {8'h00}, /* 0x70c0 */
            {8'h00}, /* 0x70bf */
            {8'h00}, /* 0x70be */
            {8'h00}, /* 0x70bd */
            {8'h00}, /* 0x70bc */
            {8'h00}, /* 0x70bb */
            {8'h00}, /* 0x70ba */
            {8'h00}, /* 0x70b9 */
            {8'h00}, /* 0x70b8 */
            {8'h00}, /* 0x70b7 */
            {8'h00}, /* 0x70b6 */
            {8'h00}, /* 0x70b5 */
            {8'h00}, /* 0x70b4 */
            {8'h00}, /* 0x70b3 */
            {8'h00}, /* 0x70b2 */
            {8'h00}, /* 0x70b1 */
            {8'h00}, /* 0x70b0 */
            {8'h00}, /* 0x70af */
            {8'h00}, /* 0x70ae */
            {8'h00}, /* 0x70ad */
            {8'h00}, /* 0x70ac */
            {8'h00}, /* 0x70ab */
            {8'h00}, /* 0x70aa */
            {8'h00}, /* 0x70a9 */
            {8'h00}, /* 0x70a8 */
            {8'h00}, /* 0x70a7 */
            {8'h00}, /* 0x70a6 */
            {8'h00}, /* 0x70a5 */
            {8'h00}, /* 0x70a4 */
            {8'h00}, /* 0x70a3 */
            {8'h00}, /* 0x70a2 */
            {8'h00}, /* 0x70a1 */
            {8'h00}, /* 0x70a0 */
            {8'h00}, /* 0x709f */
            {8'h00}, /* 0x709e */
            {8'h00}, /* 0x709d */
            {8'h00}, /* 0x709c */
            {8'h00}, /* 0x709b */
            {8'h00}, /* 0x709a */
            {8'h00}, /* 0x7099 */
            {8'h00}, /* 0x7098 */
            {8'h00}, /* 0x7097 */
            {8'h00}, /* 0x7096 */
            {8'h00}, /* 0x7095 */
            {8'h00}, /* 0x7094 */
            {8'h00}, /* 0x7093 */
            {8'h00}, /* 0x7092 */
            {8'h00}, /* 0x7091 */
            {8'h00}, /* 0x7090 */
            {8'h00}, /* 0x708f */
            {8'h00}, /* 0x708e */
            {8'h00}, /* 0x708d */
            {8'h00}, /* 0x708c */
            {8'h00}, /* 0x708b */
            {8'h00}, /* 0x708a */
            {8'h00}, /* 0x7089 */
            {8'h00}, /* 0x7088 */
            {8'h00}, /* 0x7087 */
            {8'h00}, /* 0x7086 */
            {8'h00}, /* 0x7085 */
            {8'h00}, /* 0x7084 */
            {8'h00}, /* 0x7083 */
            {8'h00}, /* 0x7082 */
            {8'h00}, /* 0x7081 */
            {8'h00}, /* 0x7080 */
            {8'h00}, /* 0x707f */
            {8'h00}, /* 0x707e */
            {8'h00}, /* 0x707d */
            {8'h00}, /* 0x707c */
            {8'h00}, /* 0x707b */
            {8'h00}, /* 0x707a */
            {8'h00}, /* 0x7079 */
            {8'h00}, /* 0x7078 */
            {8'h00}, /* 0x7077 */
            {8'h00}, /* 0x7076 */
            {8'h00}, /* 0x7075 */
            {8'h00}, /* 0x7074 */
            {8'h00}, /* 0x7073 */
            {8'h00}, /* 0x7072 */
            {8'h00}, /* 0x7071 */
            {8'h00}, /* 0x7070 */
            {8'h00}, /* 0x706f */
            {8'h00}, /* 0x706e */
            {8'h00}, /* 0x706d */
            {8'h00}, /* 0x706c */
            {8'h00}, /* 0x706b */
            {8'h00}, /* 0x706a */
            {8'h00}, /* 0x7069 */
            {8'h00}, /* 0x7068 */
            {8'h00}, /* 0x7067 */
            {8'h00}, /* 0x7066 */
            {8'h00}, /* 0x7065 */
            {8'h00}, /* 0x7064 */
            {8'h00}, /* 0x7063 */
            {8'h00}, /* 0x7062 */
            {8'h00}, /* 0x7061 */
            {8'h00}, /* 0x7060 */
            {8'h00}, /* 0x705f */
            {8'h00}, /* 0x705e */
            {8'h00}, /* 0x705d */
            {8'h00}, /* 0x705c */
            {8'h00}, /* 0x705b */
            {8'h00}, /* 0x705a */
            {8'h00}, /* 0x7059 */
            {8'h00}, /* 0x7058 */
            {8'h00}, /* 0x7057 */
            {8'h00}, /* 0x7056 */
            {8'h00}, /* 0x7055 */
            {8'h00}, /* 0x7054 */
            {8'h00}, /* 0x7053 */
            {8'h00}, /* 0x7052 */
            {8'h00}, /* 0x7051 */
            {8'h00}, /* 0x7050 */
            {8'h00}, /* 0x704f */
            {8'h00}, /* 0x704e */
            {8'h00}, /* 0x704d */
            {8'h00}, /* 0x704c */
            {8'h00}, /* 0x704b */
            {8'h00}, /* 0x704a */
            {8'h00}, /* 0x7049 */
            {8'h00}, /* 0x7048 */
            {8'h00}, /* 0x7047 */
            {8'h00}, /* 0x7046 */
            {8'h00}, /* 0x7045 */
            {8'h00}, /* 0x7044 */
            {8'h00}, /* 0x7043 */
            {8'h00}, /* 0x7042 */
            {8'h00}, /* 0x7041 */
            {8'h00}, /* 0x7040 */
            {8'h00}, /* 0x703f */
            {8'h00}, /* 0x703e */
            {8'h00}, /* 0x703d */
            {8'h00}, /* 0x703c */
            {8'h00}, /* 0x703b */
            {8'h00}, /* 0x703a */
            {8'h00}, /* 0x7039 */
            {8'h00}, /* 0x7038 */
            {8'h00}, /* 0x7037 */
            {8'h00}, /* 0x7036 */
            {8'h00}, /* 0x7035 */
            {8'h00}, /* 0x7034 */
            {8'h00}, /* 0x7033 */
            {8'h00}, /* 0x7032 */
            {8'h00}, /* 0x7031 */
            {8'h00}, /* 0x7030 */
            {8'h00}, /* 0x702f */
            {8'h00}, /* 0x702e */
            {8'h00}, /* 0x702d */
            {8'h00}, /* 0x702c */
            {8'h00}, /* 0x702b */
            {8'h00}, /* 0x702a */
            {8'h00}, /* 0x7029 */
            {8'h00}, /* 0x7028 */
            {8'h00}, /* 0x7027 */
            {8'h00}, /* 0x7026 */
            {8'h00}, /* 0x7025 */
            {8'h00}, /* 0x7024 */
            {8'h00}, /* 0x7023 */
            {8'h00}, /* 0x7022 */
            {8'h00}, /* 0x7021 */
            {8'h00}, /* 0x7020 */
            {8'h00}, /* 0x701f */
            {8'h00}, /* 0x701e */
            {8'h00}, /* 0x701d */
            {8'h00}, /* 0x701c */
            {8'h00}, /* 0x701b */
            {8'h00}, /* 0x701a */
            {8'h00}, /* 0x7019 */
            {8'h00}, /* 0x7018 */
            {8'h00}, /* 0x7017 */
            {8'h00}, /* 0x7016 */
            {8'h00}, /* 0x7015 */
            {8'h00}, /* 0x7014 */
            {8'h00}, /* 0x7013 */
            {8'h00}, /* 0x7012 */
            {8'h00}, /* 0x7011 */
            {8'h00}, /* 0x7010 */
            {8'h00}, /* 0x700f */
            {8'h00}, /* 0x700e */
            {8'h00}, /* 0x700d */
            {8'h00}, /* 0x700c */
            {8'h00}, /* 0x700b */
            {8'h00}, /* 0x700a */
            {8'h00}, /* 0x7009 */
            {8'h00}, /* 0x7008 */
            {8'h00}, /* 0x7007 */
            {8'h00}, /* 0x7006 */
            {8'h00}, /* 0x7005 */
            {8'h00}, /* 0x7004 */
            {8'h00}, /* 0x7003 */
            {8'h00}, /* 0x7002 */
            {8'h00}, /* 0x7001 */
            {8'h00}, /* 0x7000 */
            {8'h00}, /* 0x6fff */
            {8'h00}, /* 0x6ffe */
            {8'h00}, /* 0x6ffd */
            {8'h00}, /* 0x6ffc */
            {8'h00}, /* 0x6ffb */
            {8'h00}, /* 0x6ffa */
            {8'h00}, /* 0x6ff9 */
            {8'h00}, /* 0x6ff8 */
            {8'h00}, /* 0x6ff7 */
            {8'h00}, /* 0x6ff6 */
            {8'h00}, /* 0x6ff5 */
            {8'h00}, /* 0x6ff4 */
            {8'h00}, /* 0x6ff3 */
            {8'h00}, /* 0x6ff2 */
            {8'h00}, /* 0x6ff1 */
            {8'h00}, /* 0x6ff0 */
            {8'h00}, /* 0x6fef */
            {8'h00}, /* 0x6fee */
            {8'h00}, /* 0x6fed */
            {8'h00}, /* 0x6fec */
            {8'h00}, /* 0x6feb */
            {8'h00}, /* 0x6fea */
            {8'h00}, /* 0x6fe9 */
            {8'h00}, /* 0x6fe8 */
            {8'h00}, /* 0x6fe7 */
            {8'h00}, /* 0x6fe6 */
            {8'h00}, /* 0x6fe5 */
            {8'h00}, /* 0x6fe4 */
            {8'h00}, /* 0x6fe3 */
            {8'h00}, /* 0x6fe2 */
            {8'h00}, /* 0x6fe1 */
            {8'h00}, /* 0x6fe0 */
            {8'h00}, /* 0x6fdf */
            {8'h00}, /* 0x6fde */
            {8'h00}, /* 0x6fdd */
            {8'h00}, /* 0x6fdc */
            {8'h00}, /* 0x6fdb */
            {8'h00}, /* 0x6fda */
            {8'h00}, /* 0x6fd9 */
            {8'h00}, /* 0x6fd8 */
            {8'h00}, /* 0x6fd7 */
            {8'h00}, /* 0x6fd6 */
            {8'h00}, /* 0x6fd5 */
            {8'h00}, /* 0x6fd4 */
            {8'h00}, /* 0x6fd3 */
            {8'h00}, /* 0x6fd2 */
            {8'h00}, /* 0x6fd1 */
            {8'h00}, /* 0x6fd0 */
            {8'h00}, /* 0x6fcf */
            {8'h00}, /* 0x6fce */
            {8'h00}, /* 0x6fcd */
            {8'h00}, /* 0x6fcc */
            {8'h00}, /* 0x6fcb */
            {8'h00}, /* 0x6fca */
            {8'h00}, /* 0x6fc9 */
            {8'h00}, /* 0x6fc8 */
            {8'h00}, /* 0x6fc7 */
            {8'h00}, /* 0x6fc6 */
            {8'h00}, /* 0x6fc5 */
            {8'h00}, /* 0x6fc4 */
            {8'h00}, /* 0x6fc3 */
            {8'h00}, /* 0x6fc2 */
            {8'h00}, /* 0x6fc1 */
            {8'h00}, /* 0x6fc0 */
            {8'h00}, /* 0x6fbf */
            {8'h00}, /* 0x6fbe */
            {8'h00}, /* 0x6fbd */
            {8'h00}, /* 0x6fbc */
            {8'h00}, /* 0x6fbb */
            {8'h00}, /* 0x6fba */
            {8'h00}, /* 0x6fb9 */
            {8'h00}, /* 0x6fb8 */
            {8'h00}, /* 0x6fb7 */
            {8'h00}, /* 0x6fb6 */
            {8'h00}, /* 0x6fb5 */
            {8'h00}, /* 0x6fb4 */
            {8'h00}, /* 0x6fb3 */
            {8'h00}, /* 0x6fb2 */
            {8'h00}, /* 0x6fb1 */
            {8'h00}, /* 0x6fb0 */
            {8'h00}, /* 0x6faf */
            {8'h00}, /* 0x6fae */
            {8'h00}, /* 0x6fad */
            {8'h00}, /* 0x6fac */
            {8'h00}, /* 0x6fab */
            {8'h00}, /* 0x6faa */
            {8'h00}, /* 0x6fa9 */
            {8'h00}, /* 0x6fa8 */
            {8'h00}, /* 0x6fa7 */
            {8'h00}, /* 0x6fa6 */
            {8'h00}, /* 0x6fa5 */
            {8'h00}, /* 0x6fa4 */
            {8'h00}, /* 0x6fa3 */
            {8'h00}, /* 0x6fa2 */
            {8'h00}, /* 0x6fa1 */
            {8'h00}, /* 0x6fa0 */
            {8'h00}, /* 0x6f9f */
            {8'h00}, /* 0x6f9e */
            {8'h00}, /* 0x6f9d */
            {8'h00}, /* 0x6f9c */
            {8'h00}, /* 0x6f9b */
            {8'h00}, /* 0x6f9a */
            {8'h00}, /* 0x6f99 */
            {8'h00}, /* 0x6f98 */
            {8'h00}, /* 0x6f97 */
            {8'h00}, /* 0x6f96 */
            {8'h00}, /* 0x6f95 */
            {8'h00}, /* 0x6f94 */
            {8'h00}, /* 0x6f93 */
            {8'h00}, /* 0x6f92 */
            {8'h00}, /* 0x6f91 */
            {8'h00}, /* 0x6f90 */
            {8'h00}, /* 0x6f8f */
            {8'h00}, /* 0x6f8e */
            {8'h00}, /* 0x6f8d */
            {8'h00}, /* 0x6f8c */
            {8'h00}, /* 0x6f8b */
            {8'h00}, /* 0x6f8a */
            {8'h00}, /* 0x6f89 */
            {8'h00}, /* 0x6f88 */
            {8'h00}, /* 0x6f87 */
            {8'h00}, /* 0x6f86 */
            {8'h00}, /* 0x6f85 */
            {8'h00}, /* 0x6f84 */
            {8'h00}, /* 0x6f83 */
            {8'h00}, /* 0x6f82 */
            {8'h00}, /* 0x6f81 */
            {8'h00}, /* 0x6f80 */
            {8'h00}, /* 0x6f7f */
            {8'h00}, /* 0x6f7e */
            {8'h00}, /* 0x6f7d */
            {8'h00}, /* 0x6f7c */
            {8'h00}, /* 0x6f7b */
            {8'h00}, /* 0x6f7a */
            {8'h00}, /* 0x6f79 */
            {8'h00}, /* 0x6f78 */
            {8'h00}, /* 0x6f77 */
            {8'h00}, /* 0x6f76 */
            {8'h00}, /* 0x6f75 */
            {8'h00}, /* 0x6f74 */
            {8'h00}, /* 0x6f73 */
            {8'h00}, /* 0x6f72 */
            {8'h00}, /* 0x6f71 */
            {8'h00}, /* 0x6f70 */
            {8'h00}, /* 0x6f6f */
            {8'h00}, /* 0x6f6e */
            {8'h00}, /* 0x6f6d */
            {8'h00}, /* 0x6f6c */
            {8'h00}, /* 0x6f6b */
            {8'h00}, /* 0x6f6a */
            {8'h00}, /* 0x6f69 */
            {8'h00}, /* 0x6f68 */
            {8'h00}, /* 0x6f67 */
            {8'h00}, /* 0x6f66 */
            {8'h00}, /* 0x6f65 */
            {8'h00}, /* 0x6f64 */
            {8'h00}, /* 0x6f63 */
            {8'h00}, /* 0x6f62 */
            {8'h00}, /* 0x6f61 */
            {8'h00}, /* 0x6f60 */
            {8'h00}, /* 0x6f5f */
            {8'h00}, /* 0x6f5e */
            {8'h00}, /* 0x6f5d */
            {8'h00}, /* 0x6f5c */
            {8'h00}, /* 0x6f5b */
            {8'h00}, /* 0x6f5a */
            {8'h00}, /* 0x6f59 */
            {8'h00}, /* 0x6f58 */
            {8'h00}, /* 0x6f57 */
            {8'h00}, /* 0x6f56 */
            {8'h00}, /* 0x6f55 */
            {8'h00}, /* 0x6f54 */
            {8'h00}, /* 0x6f53 */
            {8'h00}, /* 0x6f52 */
            {8'h00}, /* 0x6f51 */
            {8'h00}, /* 0x6f50 */
            {8'h00}, /* 0x6f4f */
            {8'h00}, /* 0x6f4e */
            {8'h00}, /* 0x6f4d */
            {8'h00}, /* 0x6f4c */
            {8'h00}, /* 0x6f4b */
            {8'h00}, /* 0x6f4a */
            {8'h00}, /* 0x6f49 */
            {8'h00}, /* 0x6f48 */
            {8'h00}, /* 0x6f47 */
            {8'h00}, /* 0x6f46 */
            {8'h00}, /* 0x6f45 */
            {8'h00}, /* 0x6f44 */
            {8'h00}, /* 0x6f43 */
            {8'h00}, /* 0x6f42 */
            {8'h00}, /* 0x6f41 */
            {8'h00}, /* 0x6f40 */
            {8'h00}, /* 0x6f3f */
            {8'h00}, /* 0x6f3e */
            {8'h00}, /* 0x6f3d */
            {8'h00}, /* 0x6f3c */
            {8'h00}, /* 0x6f3b */
            {8'h00}, /* 0x6f3a */
            {8'h00}, /* 0x6f39 */
            {8'h00}, /* 0x6f38 */
            {8'h00}, /* 0x6f37 */
            {8'h00}, /* 0x6f36 */
            {8'h00}, /* 0x6f35 */
            {8'h00}, /* 0x6f34 */
            {8'h00}, /* 0x6f33 */
            {8'h00}, /* 0x6f32 */
            {8'h00}, /* 0x6f31 */
            {8'h00}, /* 0x6f30 */
            {8'h00}, /* 0x6f2f */
            {8'h00}, /* 0x6f2e */
            {8'h00}, /* 0x6f2d */
            {8'h00}, /* 0x6f2c */
            {8'h00}, /* 0x6f2b */
            {8'h00}, /* 0x6f2a */
            {8'h00}, /* 0x6f29 */
            {8'h00}, /* 0x6f28 */
            {8'h00}, /* 0x6f27 */
            {8'h00}, /* 0x6f26 */
            {8'h00}, /* 0x6f25 */
            {8'h00}, /* 0x6f24 */
            {8'h00}, /* 0x6f23 */
            {8'h00}, /* 0x6f22 */
            {8'h00}, /* 0x6f21 */
            {8'h00}, /* 0x6f20 */
            {8'h00}, /* 0x6f1f */
            {8'h00}, /* 0x6f1e */
            {8'h00}, /* 0x6f1d */
            {8'h00}, /* 0x6f1c */
            {8'h00}, /* 0x6f1b */
            {8'h00}, /* 0x6f1a */
            {8'h00}, /* 0x6f19 */
            {8'h00}, /* 0x6f18 */
            {8'h00}, /* 0x6f17 */
            {8'h00}, /* 0x6f16 */
            {8'h00}, /* 0x6f15 */
            {8'h00}, /* 0x6f14 */
            {8'h00}, /* 0x6f13 */
            {8'h00}, /* 0x6f12 */
            {8'h00}, /* 0x6f11 */
            {8'h00}, /* 0x6f10 */
            {8'h00}, /* 0x6f0f */
            {8'h00}, /* 0x6f0e */
            {8'h00}, /* 0x6f0d */
            {8'h00}, /* 0x6f0c */
            {8'h00}, /* 0x6f0b */
            {8'h00}, /* 0x6f0a */
            {8'h00}, /* 0x6f09 */
            {8'h00}, /* 0x6f08 */
            {8'h00}, /* 0x6f07 */
            {8'h00}, /* 0x6f06 */
            {8'h00}, /* 0x6f05 */
            {8'h00}, /* 0x6f04 */
            {8'h00}, /* 0x6f03 */
            {8'h00}, /* 0x6f02 */
            {8'h00}, /* 0x6f01 */
            {8'h00}, /* 0x6f00 */
            {8'h00}, /* 0x6eff */
            {8'h00}, /* 0x6efe */
            {8'h00}, /* 0x6efd */
            {8'h00}, /* 0x6efc */
            {8'h00}, /* 0x6efb */
            {8'h00}, /* 0x6efa */
            {8'h00}, /* 0x6ef9 */
            {8'h00}, /* 0x6ef8 */
            {8'h00}, /* 0x6ef7 */
            {8'h00}, /* 0x6ef6 */
            {8'h00}, /* 0x6ef5 */
            {8'h00}, /* 0x6ef4 */
            {8'h00}, /* 0x6ef3 */
            {8'h00}, /* 0x6ef2 */
            {8'h00}, /* 0x6ef1 */
            {8'h00}, /* 0x6ef0 */
            {8'h00}, /* 0x6eef */
            {8'h00}, /* 0x6eee */
            {8'h00}, /* 0x6eed */
            {8'h00}, /* 0x6eec */
            {8'h00}, /* 0x6eeb */
            {8'h00}, /* 0x6eea */
            {8'h00}, /* 0x6ee9 */
            {8'h00}, /* 0x6ee8 */
            {8'h00}, /* 0x6ee7 */
            {8'h00}, /* 0x6ee6 */
            {8'h00}, /* 0x6ee5 */
            {8'h00}, /* 0x6ee4 */
            {8'h00}, /* 0x6ee3 */
            {8'h00}, /* 0x6ee2 */
            {8'h00}, /* 0x6ee1 */
            {8'h00}, /* 0x6ee0 */
            {8'h00}, /* 0x6edf */
            {8'h00}, /* 0x6ede */
            {8'h00}, /* 0x6edd */
            {8'h00}, /* 0x6edc */
            {8'h00}, /* 0x6edb */
            {8'h00}, /* 0x6eda */
            {8'h00}, /* 0x6ed9 */
            {8'h00}, /* 0x6ed8 */
            {8'h00}, /* 0x6ed7 */
            {8'h00}, /* 0x6ed6 */
            {8'h00}, /* 0x6ed5 */
            {8'h00}, /* 0x6ed4 */
            {8'h00}, /* 0x6ed3 */
            {8'h00}, /* 0x6ed2 */
            {8'h00}, /* 0x6ed1 */
            {8'h00}, /* 0x6ed0 */
            {8'h00}, /* 0x6ecf */
            {8'h00}, /* 0x6ece */
            {8'h00}, /* 0x6ecd */
            {8'h00}, /* 0x6ecc */
            {8'h00}, /* 0x6ecb */
            {8'h00}, /* 0x6eca */
            {8'h00}, /* 0x6ec9 */
            {8'h00}, /* 0x6ec8 */
            {8'h00}, /* 0x6ec7 */
            {8'h00}, /* 0x6ec6 */
            {8'h00}, /* 0x6ec5 */
            {8'h00}, /* 0x6ec4 */
            {8'h00}, /* 0x6ec3 */
            {8'h00}, /* 0x6ec2 */
            {8'h00}, /* 0x6ec1 */
            {8'h00}, /* 0x6ec0 */
            {8'h00}, /* 0x6ebf */
            {8'h00}, /* 0x6ebe */
            {8'h00}, /* 0x6ebd */
            {8'h00}, /* 0x6ebc */
            {8'h00}, /* 0x6ebb */
            {8'h00}, /* 0x6eba */
            {8'h00}, /* 0x6eb9 */
            {8'h00}, /* 0x6eb8 */
            {8'h00}, /* 0x6eb7 */
            {8'h00}, /* 0x6eb6 */
            {8'h00}, /* 0x6eb5 */
            {8'h00}, /* 0x6eb4 */
            {8'h00}, /* 0x6eb3 */
            {8'h00}, /* 0x6eb2 */
            {8'h00}, /* 0x6eb1 */
            {8'h00}, /* 0x6eb0 */
            {8'h00}, /* 0x6eaf */
            {8'h00}, /* 0x6eae */
            {8'h00}, /* 0x6ead */
            {8'h00}, /* 0x6eac */
            {8'h00}, /* 0x6eab */
            {8'h00}, /* 0x6eaa */
            {8'h00}, /* 0x6ea9 */
            {8'h00}, /* 0x6ea8 */
            {8'h00}, /* 0x6ea7 */
            {8'h00}, /* 0x6ea6 */
            {8'h00}, /* 0x6ea5 */
            {8'h00}, /* 0x6ea4 */
            {8'h00}, /* 0x6ea3 */
            {8'h00}, /* 0x6ea2 */
            {8'h00}, /* 0x6ea1 */
            {8'h00}, /* 0x6ea0 */
            {8'h00}, /* 0x6e9f */
            {8'h00}, /* 0x6e9e */
            {8'h00}, /* 0x6e9d */
            {8'h00}, /* 0x6e9c */
            {8'h00}, /* 0x6e9b */
            {8'h00}, /* 0x6e9a */
            {8'h00}, /* 0x6e99 */
            {8'h00}, /* 0x6e98 */
            {8'h00}, /* 0x6e97 */
            {8'h00}, /* 0x6e96 */
            {8'h00}, /* 0x6e95 */
            {8'h00}, /* 0x6e94 */
            {8'h00}, /* 0x6e93 */
            {8'h00}, /* 0x6e92 */
            {8'h00}, /* 0x6e91 */
            {8'h00}, /* 0x6e90 */
            {8'h00}, /* 0x6e8f */
            {8'h00}, /* 0x6e8e */
            {8'h00}, /* 0x6e8d */
            {8'h00}, /* 0x6e8c */
            {8'h00}, /* 0x6e8b */
            {8'h00}, /* 0x6e8a */
            {8'h00}, /* 0x6e89 */
            {8'h00}, /* 0x6e88 */
            {8'h00}, /* 0x6e87 */
            {8'h00}, /* 0x6e86 */
            {8'h00}, /* 0x6e85 */
            {8'h00}, /* 0x6e84 */
            {8'h00}, /* 0x6e83 */
            {8'h00}, /* 0x6e82 */
            {8'h00}, /* 0x6e81 */
            {8'h00}, /* 0x6e80 */
            {8'h00}, /* 0x6e7f */
            {8'h00}, /* 0x6e7e */
            {8'h00}, /* 0x6e7d */
            {8'h00}, /* 0x6e7c */
            {8'h00}, /* 0x6e7b */
            {8'h00}, /* 0x6e7a */
            {8'h00}, /* 0x6e79 */
            {8'h00}, /* 0x6e78 */
            {8'h00}, /* 0x6e77 */
            {8'h00}, /* 0x6e76 */
            {8'h00}, /* 0x6e75 */
            {8'h00}, /* 0x6e74 */
            {8'h00}, /* 0x6e73 */
            {8'h00}, /* 0x6e72 */
            {8'h00}, /* 0x6e71 */
            {8'h00}, /* 0x6e70 */
            {8'h00}, /* 0x6e6f */
            {8'h00}, /* 0x6e6e */
            {8'h00}, /* 0x6e6d */
            {8'h00}, /* 0x6e6c */
            {8'h00}, /* 0x6e6b */
            {8'h00}, /* 0x6e6a */
            {8'h00}, /* 0x6e69 */
            {8'h00}, /* 0x6e68 */
            {8'h00}, /* 0x6e67 */
            {8'h00}, /* 0x6e66 */
            {8'h00}, /* 0x6e65 */
            {8'h00}, /* 0x6e64 */
            {8'h00}, /* 0x6e63 */
            {8'h00}, /* 0x6e62 */
            {8'h00}, /* 0x6e61 */
            {8'h00}, /* 0x6e60 */
            {8'h00}, /* 0x6e5f */
            {8'h00}, /* 0x6e5e */
            {8'h00}, /* 0x6e5d */
            {8'h00}, /* 0x6e5c */
            {8'h00}, /* 0x6e5b */
            {8'h00}, /* 0x6e5a */
            {8'h00}, /* 0x6e59 */
            {8'h00}, /* 0x6e58 */
            {8'h00}, /* 0x6e57 */
            {8'h00}, /* 0x6e56 */
            {8'h00}, /* 0x6e55 */
            {8'h00}, /* 0x6e54 */
            {8'h00}, /* 0x6e53 */
            {8'h00}, /* 0x6e52 */
            {8'h00}, /* 0x6e51 */
            {8'h00}, /* 0x6e50 */
            {8'h00}, /* 0x6e4f */
            {8'h00}, /* 0x6e4e */
            {8'h00}, /* 0x6e4d */
            {8'h00}, /* 0x6e4c */
            {8'h00}, /* 0x6e4b */
            {8'h00}, /* 0x6e4a */
            {8'h00}, /* 0x6e49 */
            {8'h00}, /* 0x6e48 */
            {8'h00}, /* 0x6e47 */
            {8'h00}, /* 0x6e46 */
            {8'h00}, /* 0x6e45 */
            {8'h00}, /* 0x6e44 */
            {8'h00}, /* 0x6e43 */
            {8'h00}, /* 0x6e42 */
            {8'h00}, /* 0x6e41 */
            {8'h00}, /* 0x6e40 */
            {8'h00}, /* 0x6e3f */
            {8'h00}, /* 0x6e3e */
            {8'h00}, /* 0x6e3d */
            {8'h00}, /* 0x6e3c */
            {8'h00}, /* 0x6e3b */
            {8'h00}, /* 0x6e3a */
            {8'h00}, /* 0x6e39 */
            {8'h00}, /* 0x6e38 */
            {8'h00}, /* 0x6e37 */
            {8'h00}, /* 0x6e36 */
            {8'h00}, /* 0x6e35 */
            {8'h00}, /* 0x6e34 */
            {8'h00}, /* 0x6e33 */
            {8'h00}, /* 0x6e32 */
            {8'h00}, /* 0x6e31 */
            {8'h00}, /* 0x6e30 */
            {8'h00}, /* 0x6e2f */
            {8'h00}, /* 0x6e2e */
            {8'h00}, /* 0x6e2d */
            {8'h00}, /* 0x6e2c */
            {8'h00}, /* 0x6e2b */
            {8'h00}, /* 0x6e2a */
            {8'h00}, /* 0x6e29 */
            {8'h00}, /* 0x6e28 */
            {8'h00}, /* 0x6e27 */
            {8'h00}, /* 0x6e26 */
            {8'h00}, /* 0x6e25 */
            {8'h00}, /* 0x6e24 */
            {8'h00}, /* 0x6e23 */
            {8'h00}, /* 0x6e22 */
            {8'h00}, /* 0x6e21 */
            {8'h00}, /* 0x6e20 */
            {8'h00}, /* 0x6e1f */
            {8'h00}, /* 0x6e1e */
            {8'h00}, /* 0x6e1d */
            {8'h00}, /* 0x6e1c */
            {8'h00}, /* 0x6e1b */
            {8'h00}, /* 0x6e1a */
            {8'h00}, /* 0x6e19 */
            {8'h00}, /* 0x6e18 */
            {8'h00}, /* 0x6e17 */
            {8'h00}, /* 0x6e16 */
            {8'h00}, /* 0x6e15 */
            {8'h00}, /* 0x6e14 */
            {8'h00}, /* 0x6e13 */
            {8'h00}, /* 0x6e12 */
            {8'h00}, /* 0x6e11 */
            {8'h00}, /* 0x6e10 */
            {8'h00}, /* 0x6e0f */
            {8'h00}, /* 0x6e0e */
            {8'h00}, /* 0x6e0d */
            {8'h00}, /* 0x6e0c */
            {8'h00}, /* 0x6e0b */
            {8'h00}, /* 0x6e0a */
            {8'h00}, /* 0x6e09 */
            {8'h00}, /* 0x6e08 */
            {8'h00}, /* 0x6e07 */
            {8'h00}, /* 0x6e06 */
            {8'h00}, /* 0x6e05 */
            {8'h00}, /* 0x6e04 */
            {8'h00}, /* 0x6e03 */
            {8'h00}, /* 0x6e02 */
            {8'h00}, /* 0x6e01 */
            {8'h00}, /* 0x6e00 */
            {8'h00}, /* 0x6dff */
            {8'h00}, /* 0x6dfe */
            {8'h00}, /* 0x6dfd */
            {8'h00}, /* 0x6dfc */
            {8'h00}, /* 0x6dfb */
            {8'h00}, /* 0x6dfa */
            {8'h00}, /* 0x6df9 */
            {8'h00}, /* 0x6df8 */
            {8'h00}, /* 0x6df7 */
            {8'h00}, /* 0x6df6 */
            {8'h00}, /* 0x6df5 */
            {8'h00}, /* 0x6df4 */
            {8'h00}, /* 0x6df3 */
            {8'h00}, /* 0x6df2 */
            {8'h00}, /* 0x6df1 */
            {8'h00}, /* 0x6df0 */
            {8'h00}, /* 0x6def */
            {8'h00}, /* 0x6dee */
            {8'h00}, /* 0x6ded */
            {8'h00}, /* 0x6dec */
            {8'h00}, /* 0x6deb */
            {8'h00}, /* 0x6dea */
            {8'h00}, /* 0x6de9 */
            {8'h00}, /* 0x6de8 */
            {8'h00}, /* 0x6de7 */
            {8'h00}, /* 0x6de6 */
            {8'h00}, /* 0x6de5 */
            {8'h00}, /* 0x6de4 */
            {8'h00}, /* 0x6de3 */
            {8'h00}, /* 0x6de2 */
            {8'h00}, /* 0x6de1 */
            {8'h00}, /* 0x6de0 */
            {8'h00}, /* 0x6ddf */
            {8'h00}, /* 0x6dde */
            {8'h00}, /* 0x6ddd */
            {8'h00}, /* 0x6ddc */
            {8'h00}, /* 0x6ddb */
            {8'h00}, /* 0x6dda */
            {8'h00}, /* 0x6dd9 */
            {8'h00}, /* 0x6dd8 */
            {8'h00}, /* 0x6dd7 */
            {8'h00}, /* 0x6dd6 */
            {8'h00}, /* 0x6dd5 */
            {8'h00}, /* 0x6dd4 */
            {8'h00}, /* 0x6dd3 */
            {8'h00}, /* 0x6dd2 */
            {8'h00}, /* 0x6dd1 */
            {8'h00}, /* 0x6dd0 */
            {8'h00}, /* 0x6dcf */
            {8'h00}, /* 0x6dce */
            {8'h00}, /* 0x6dcd */
            {8'h00}, /* 0x6dcc */
            {8'h00}, /* 0x6dcb */
            {8'h00}, /* 0x6dca */
            {8'h00}, /* 0x6dc9 */
            {8'h00}, /* 0x6dc8 */
            {8'h00}, /* 0x6dc7 */
            {8'h00}, /* 0x6dc6 */
            {8'h00}, /* 0x6dc5 */
            {8'h00}, /* 0x6dc4 */
            {8'h00}, /* 0x6dc3 */
            {8'h00}, /* 0x6dc2 */
            {8'h00}, /* 0x6dc1 */
            {8'h00}, /* 0x6dc0 */
            {8'h00}, /* 0x6dbf */
            {8'h00}, /* 0x6dbe */
            {8'h00}, /* 0x6dbd */
            {8'h00}, /* 0x6dbc */
            {8'h00}, /* 0x6dbb */
            {8'h00}, /* 0x6dba */
            {8'h00}, /* 0x6db9 */
            {8'h00}, /* 0x6db8 */
            {8'h00}, /* 0x6db7 */
            {8'h00}, /* 0x6db6 */
            {8'h00}, /* 0x6db5 */
            {8'h00}, /* 0x6db4 */
            {8'h00}, /* 0x6db3 */
            {8'h00}, /* 0x6db2 */
            {8'h00}, /* 0x6db1 */
            {8'h00}, /* 0x6db0 */
            {8'h00}, /* 0x6daf */
            {8'h00}, /* 0x6dae */
            {8'h00}, /* 0x6dad */
            {8'h00}, /* 0x6dac */
            {8'h00}, /* 0x6dab */
            {8'h00}, /* 0x6daa */
            {8'h00}, /* 0x6da9 */
            {8'h00}, /* 0x6da8 */
            {8'h00}, /* 0x6da7 */
            {8'h00}, /* 0x6da6 */
            {8'h00}, /* 0x6da5 */
            {8'h00}, /* 0x6da4 */
            {8'h00}, /* 0x6da3 */
            {8'h00}, /* 0x6da2 */
            {8'h00}, /* 0x6da1 */
            {8'h00}, /* 0x6da0 */
            {8'h00}, /* 0x6d9f */
            {8'h00}, /* 0x6d9e */
            {8'h00}, /* 0x6d9d */
            {8'h00}, /* 0x6d9c */
            {8'h00}, /* 0x6d9b */
            {8'h00}, /* 0x6d9a */
            {8'h00}, /* 0x6d99 */
            {8'h00}, /* 0x6d98 */
            {8'h00}, /* 0x6d97 */
            {8'h00}, /* 0x6d96 */
            {8'h00}, /* 0x6d95 */
            {8'h00}, /* 0x6d94 */
            {8'h00}, /* 0x6d93 */
            {8'h00}, /* 0x6d92 */
            {8'h00}, /* 0x6d91 */
            {8'h00}, /* 0x6d90 */
            {8'h00}, /* 0x6d8f */
            {8'h00}, /* 0x6d8e */
            {8'h00}, /* 0x6d8d */
            {8'h00}, /* 0x6d8c */
            {8'h00}, /* 0x6d8b */
            {8'h00}, /* 0x6d8a */
            {8'h00}, /* 0x6d89 */
            {8'h00}, /* 0x6d88 */
            {8'h00}, /* 0x6d87 */
            {8'h00}, /* 0x6d86 */
            {8'h00}, /* 0x6d85 */
            {8'h00}, /* 0x6d84 */
            {8'h00}, /* 0x6d83 */
            {8'h00}, /* 0x6d82 */
            {8'h00}, /* 0x6d81 */
            {8'h00}, /* 0x6d80 */
            {8'h00}, /* 0x6d7f */
            {8'h00}, /* 0x6d7e */
            {8'h00}, /* 0x6d7d */
            {8'h00}, /* 0x6d7c */
            {8'h00}, /* 0x6d7b */
            {8'h00}, /* 0x6d7a */
            {8'h00}, /* 0x6d79 */
            {8'h00}, /* 0x6d78 */
            {8'h00}, /* 0x6d77 */
            {8'h00}, /* 0x6d76 */
            {8'h00}, /* 0x6d75 */
            {8'h00}, /* 0x6d74 */
            {8'h00}, /* 0x6d73 */
            {8'h00}, /* 0x6d72 */
            {8'h00}, /* 0x6d71 */
            {8'h00}, /* 0x6d70 */
            {8'h00}, /* 0x6d6f */
            {8'h00}, /* 0x6d6e */
            {8'h00}, /* 0x6d6d */
            {8'h00}, /* 0x6d6c */
            {8'h00}, /* 0x6d6b */
            {8'h00}, /* 0x6d6a */
            {8'h00}, /* 0x6d69 */
            {8'h00}, /* 0x6d68 */
            {8'h00}, /* 0x6d67 */
            {8'h00}, /* 0x6d66 */
            {8'h00}, /* 0x6d65 */
            {8'h00}, /* 0x6d64 */
            {8'h00}, /* 0x6d63 */
            {8'h00}, /* 0x6d62 */
            {8'h00}, /* 0x6d61 */
            {8'h00}, /* 0x6d60 */
            {8'h00}, /* 0x6d5f */
            {8'h00}, /* 0x6d5e */
            {8'h00}, /* 0x6d5d */
            {8'h00}, /* 0x6d5c */
            {8'h00}, /* 0x6d5b */
            {8'h00}, /* 0x6d5a */
            {8'h00}, /* 0x6d59 */
            {8'h00}, /* 0x6d58 */
            {8'h00}, /* 0x6d57 */
            {8'h00}, /* 0x6d56 */
            {8'h00}, /* 0x6d55 */
            {8'h00}, /* 0x6d54 */
            {8'h00}, /* 0x6d53 */
            {8'h00}, /* 0x6d52 */
            {8'h00}, /* 0x6d51 */
            {8'h00}, /* 0x6d50 */
            {8'h00}, /* 0x6d4f */
            {8'h00}, /* 0x6d4e */
            {8'h00}, /* 0x6d4d */
            {8'h00}, /* 0x6d4c */
            {8'h00}, /* 0x6d4b */
            {8'h00}, /* 0x6d4a */
            {8'h00}, /* 0x6d49 */
            {8'h00}, /* 0x6d48 */
            {8'h00}, /* 0x6d47 */
            {8'h00}, /* 0x6d46 */
            {8'h00}, /* 0x6d45 */
            {8'h00}, /* 0x6d44 */
            {8'h00}, /* 0x6d43 */
            {8'h00}, /* 0x6d42 */
            {8'h00}, /* 0x6d41 */
            {8'h00}, /* 0x6d40 */
            {8'h00}, /* 0x6d3f */
            {8'h00}, /* 0x6d3e */
            {8'h00}, /* 0x6d3d */
            {8'h00}, /* 0x6d3c */
            {8'h00}, /* 0x6d3b */
            {8'h00}, /* 0x6d3a */
            {8'h00}, /* 0x6d39 */
            {8'h00}, /* 0x6d38 */
            {8'h00}, /* 0x6d37 */
            {8'h00}, /* 0x6d36 */
            {8'h00}, /* 0x6d35 */
            {8'h00}, /* 0x6d34 */
            {8'h00}, /* 0x6d33 */
            {8'h00}, /* 0x6d32 */
            {8'h00}, /* 0x6d31 */
            {8'h00}, /* 0x6d30 */
            {8'h00}, /* 0x6d2f */
            {8'h00}, /* 0x6d2e */
            {8'h00}, /* 0x6d2d */
            {8'h00}, /* 0x6d2c */
            {8'h00}, /* 0x6d2b */
            {8'h00}, /* 0x6d2a */
            {8'h00}, /* 0x6d29 */
            {8'h00}, /* 0x6d28 */
            {8'h00}, /* 0x6d27 */
            {8'h00}, /* 0x6d26 */
            {8'h00}, /* 0x6d25 */
            {8'h00}, /* 0x6d24 */
            {8'h00}, /* 0x6d23 */
            {8'h00}, /* 0x6d22 */
            {8'h00}, /* 0x6d21 */
            {8'h00}, /* 0x6d20 */
            {8'h00}, /* 0x6d1f */
            {8'h00}, /* 0x6d1e */
            {8'h00}, /* 0x6d1d */
            {8'h00}, /* 0x6d1c */
            {8'h00}, /* 0x6d1b */
            {8'h00}, /* 0x6d1a */
            {8'h00}, /* 0x6d19 */
            {8'h00}, /* 0x6d18 */
            {8'h00}, /* 0x6d17 */
            {8'h00}, /* 0x6d16 */
            {8'h00}, /* 0x6d15 */
            {8'h00}, /* 0x6d14 */
            {8'h00}, /* 0x6d13 */
            {8'h00}, /* 0x6d12 */
            {8'h00}, /* 0x6d11 */
            {8'h00}, /* 0x6d10 */
            {8'h00}, /* 0x6d0f */
            {8'h00}, /* 0x6d0e */
            {8'h00}, /* 0x6d0d */
            {8'h00}, /* 0x6d0c */
            {8'h00}, /* 0x6d0b */
            {8'h00}, /* 0x6d0a */
            {8'h00}, /* 0x6d09 */
            {8'h00}, /* 0x6d08 */
            {8'h00}, /* 0x6d07 */
            {8'h00}, /* 0x6d06 */
            {8'h00}, /* 0x6d05 */
            {8'h00}, /* 0x6d04 */
            {8'h00}, /* 0x6d03 */
            {8'h00}, /* 0x6d02 */
            {8'h00}, /* 0x6d01 */
            {8'h00}, /* 0x6d00 */
            {8'h00}, /* 0x6cff */
            {8'h00}, /* 0x6cfe */
            {8'h00}, /* 0x6cfd */
            {8'h00}, /* 0x6cfc */
            {8'h00}, /* 0x6cfb */
            {8'h00}, /* 0x6cfa */
            {8'h00}, /* 0x6cf9 */
            {8'h00}, /* 0x6cf8 */
            {8'h00}, /* 0x6cf7 */
            {8'h00}, /* 0x6cf6 */
            {8'h00}, /* 0x6cf5 */
            {8'h00}, /* 0x6cf4 */
            {8'h00}, /* 0x6cf3 */
            {8'h00}, /* 0x6cf2 */
            {8'h00}, /* 0x6cf1 */
            {8'h00}, /* 0x6cf0 */
            {8'h00}, /* 0x6cef */
            {8'h00}, /* 0x6cee */
            {8'h00}, /* 0x6ced */
            {8'h00}, /* 0x6cec */
            {8'h00}, /* 0x6ceb */
            {8'h00}, /* 0x6cea */
            {8'h00}, /* 0x6ce9 */
            {8'h00}, /* 0x6ce8 */
            {8'h00}, /* 0x6ce7 */
            {8'h00}, /* 0x6ce6 */
            {8'h00}, /* 0x6ce5 */
            {8'h00}, /* 0x6ce4 */
            {8'h00}, /* 0x6ce3 */
            {8'h00}, /* 0x6ce2 */
            {8'h00}, /* 0x6ce1 */
            {8'h00}, /* 0x6ce0 */
            {8'h00}, /* 0x6cdf */
            {8'h00}, /* 0x6cde */
            {8'h00}, /* 0x6cdd */
            {8'h00}, /* 0x6cdc */
            {8'h00}, /* 0x6cdb */
            {8'h00}, /* 0x6cda */
            {8'h00}, /* 0x6cd9 */
            {8'h00}, /* 0x6cd8 */
            {8'h00}, /* 0x6cd7 */
            {8'h00}, /* 0x6cd6 */
            {8'h00}, /* 0x6cd5 */
            {8'h00}, /* 0x6cd4 */
            {8'h00}, /* 0x6cd3 */
            {8'h00}, /* 0x6cd2 */
            {8'h00}, /* 0x6cd1 */
            {8'h00}, /* 0x6cd0 */
            {8'h00}, /* 0x6ccf */
            {8'h00}, /* 0x6cce */
            {8'h00}, /* 0x6ccd */
            {8'h00}, /* 0x6ccc */
            {8'h00}, /* 0x6ccb */
            {8'h00}, /* 0x6cca */
            {8'h00}, /* 0x6cc9 */
            {8'h00}, /* 0x6cc8 */
            {8'h00}, /* 0x6cc7 */
            {8'h00}, /* 0x6cc6 */
            {8'h00}, /* 0x6cc5 */
            {8'h00}, /* 0x6cc4 */
            {8'h00}, /* 0x6cc3 */
            {8'h00}, /* 0x6cc2 */
            {8'h00}, /* 0x6cc1 */
            {8'h00}, /* 0x6cc0 */
            {8'h00}, /* 0x6cbf */
            {8'h00}, /* 0x6cbe */
            {8'h00}, /* 0x6cbd */
            {8'h00}, /* 0x6cbc */
            {8'h00}, /* 0x6cbb */
            {8'h00}, /* 0x6cba */
            {8'h00}, /* 0x6cb9 */
            {8'h00}, /* 0x6cb8 */
            {8'h00}, /* 0x6cb7 */
            {8'h00}, /* 0x6cb6 */
            {8'h00}, /* 0x6cb5 */
            {8'h00}, /* 0x6cb4 */
            {8'h00}, /* 0x6cb3 */
            {8'h00}, /* 0x6cb2 */
            {8'h00}, /* 0x6cb1 */
            {8'h00}, /* 0x6cb0 */
            {8'h00}, /* 0x6caf */
            {8'h00}, /* 0x6cae */
            {8'h00}, /* 0x6cad */
            {8'h00}, /* 0x6cac */
            {8'h00}, /* 0x6cab */
            {8'h00}, /* 0x6caa */
            {8'h00}, /* 0x6ca9 */
            {8'h00}, /* 0x6ca8 */
            {8'h00}, /* 0x6ca7 */
            {8'h00}, /* 0x6ca6 */
            {8'h00}, /* 0x6ca5 */
            {8'h00}, /* 0x6ca4 */
            {8'h00}, /* 0x6ca3 */
            {8'h00}, /* 0x6ca2 */
            {8'h00}, /* 0x6ca1 */
            {8'h00}, /* 0x6ca0 */
            {8'h00}, /* 0x6c9f */
            {8'h00}, /* 0x6c9e */
            {8'h00}, /* 0x6c9d */
            {8'h00}, /* 0x6c9c */
            {8'h00}, /* 0x6c9b */
            {8'h00}, /* 0x6c9a */
            {8'h00}, /* 0x6c99 */
            {8'h00}, /* 0x6c98 */
            {8'h00}, /* 0x6c97 */
            {8'h00}, /* 0x6c96 */
            {8'h00}, /* 0x6c95 */
            {8'h00}, /* 0x6c94 */
            {8'h00}, /* 0x6c93 */
            {8'h00}, /* 0x6c92 */
            {8'h00}, /* 0x6c91 */
            {8'h00}, /* 0x6c90 */
            {8'h00}, /* 0x6c8f */
            {8'h00}, /* 0x6c8e */
            {8'h00}, /* 0x6c8d */
            {8'h00}, /* 0x6c8c */
            {8'h00}, /* 0x6c8b */
            {8'h00}, /* 0x6c8a */
            {8'h00}, /* 0x6c89 */
            {8'h00}, /* 0x6c88 */
            {8'h00}, /* 0x6c87 */
            {8'h00}, /* 0x6c86 */
            {8'h00}, /* 0x6c85 */
            {8'h00}, /* 0x6c84 */
            {8'h00}, /* 0x6c83 */
            {8'h00}, /* 0x6c82 */
            {8'h00}, /* 0x6c81 */
            {8'h00}, /* 0x6c80 */
            {8'h00}, /* 0x6c7f */
            {8'h00}, /* 0x6c7e */
            {8'h00}, /* 0x6c7d */
            {8'h00}, /* 0x6c7c */
            {8'h00}, /* 0x6c7b */
            {8'h00}, /* 0x6c7a */
            {8'h00}, /* 0x6c79 */
            {8'h00}, /* 0x6c78 */
            {8'h00}, /* 0x6c77 */
            {8'h00}, /* 0x6c76 */
            {8'h00}, /* 0x6c75 */
            {8'h00}, /* 0x6c74 */
            {8'h00}, /* 0x6c73 */
            {8'h00}, /* 0x6c72 */
            {8'h00}, /* 0x6c71 */
            {8'h00}, /* 0x6c70 */
            {8'h00}, /* 0x6c6f */
            {8'h00}, /* 0x6c6e */
            {8'h00}, /* 0x6c6d */
            {8'h00}, /* 0x6c6c */
            {8'h00}, /* 0x6c6b */
            {8'h00}, /* 0x6c6a */
            {8'h00}, /* 0x6c69 */
            {8'h00}, /* 0x6c68 */
            {8'h00}, /* 0x6c67 */
            {8'h00}, /* 0x6c66 */
            {8'h00}, /* 0x6c65 */
            {8'h00}, /* 0x6c64 */
            {8'h00}, /* 0x6c63 */
            {8'h00}, /* 0x6c62 */
            {8'h00}, /* 0x6c61 */
            {8'h00}, /* 0x6c60 */
            {8'h00}, /* 0x6c5f */
            {8'h00}, /* 0x6c5e */
            {8'h00}, /* 0x6c5d */
            {8'h00}, /* 0x6c5c */
            {8'h00}, /* 0x6c5b */
            {8'h00}, /* 0x6c5a */
            {8'h00}, /* 0x6c59 */
            {8'h00}, /* 0x6c58 */
            {8'h00}, /* 0x6c57 */
            {8'h00}, /* 0x6c56 */
            {8'h00}, /* 0x6c55 */
            {8'h00}, /* 0x6c54 */
            {8'h00}, /* 0x6c53 */
            {8'h00}, /* 0x6c52 */
            {8'h00}, /* 0x6c51 */
            {8'h00}, /* 0x6c50 */
            {8'h00}, /* 0x6c4f */
            {8'h00}, /* 0x6c4e */
            {8'h00}, /* 0x6c4d */
            {8'h00}, /* 0x6c4c */
            {8'h00}, /* 0x6c4b */
            {8'h00}, /* 0x6c4a */
            {8'h00}, /* 0x6c49 */
            {8'h00}, /* 0x6c48 */
            {8'h00}, /* 0x6c47 */
            {8'h00}, /* 0x6c46 */
            {8'h00}, /* 0x6c45 */
            {8'h00}, /* 0x6c44 */
            {8'h00}, /* 0x6c43 */
            {8'h00}, /* 0x6c42 */
            {8'h00}, /* 0x6c41 */
            {8'h00}, /* 0x6c40 */
            {8'h00}, /* 0x6c3f */
            {8'h00}, /* 0x6c3e */
            {8'h00}, /* 0x6c3d */
            {8'h00}, /* 0x6c3c */
            {8'h00}, /* 0x6c3b */
            {8'h00}, /* 0x6c3a */
            {8'h00}, /* 0x6c39 */
            {8'h00}, /* 0x6c38 */
            {8'h00}, /* 0x6c37 */
            {8'h00}, /* 0x6c36 */
            {8'h00}, /* 0x6c35 */
            {8'h00}, /* 0x6c34 */
            {8'h00}, /* 0x6c33 */
            {8'h00}, /* 0x6c32 */
            {8'h00}, /* 0x6c31 */
            {8'h00}, /* 0x6c30 */
            {8'h00}, /* 0x6c2f */
            {8'h00}, /* 0x6c2e */
            {8'h00}, /* 0x6c2d */
            {8'h00}, /* 0x6c2c */
            {8'h00}, /* 0x6c2b */
            {8'h00}, /* 0x6c2a */
            {8'h00}, /* 0x6c29 */
            {8'h00}, /* 0x6c28 */
            {8'h00}, /* 0x6c27 */
            {8'h00}, /* 0x6c26 */
            {8'h00}, /* 0x6c25 */
            {8'h00}, /* 0x6c24 */
            {8'h00}, /* 0x6c23 */
            {8'h00}, /* 0x6c22 */
            {8'h00}, /* 0x6c21 */
            {8'h00}, /* 0x6c20 */
            {8'h00}, /* 0x6c1f */
            {8'h00}, /* 0x6c1e */
            {8'h00}, /* 0x6c1d */
            {8'h00}, /* 0x6c1c */
            {8'h00}, /* 0x6c1b */
            {8'h00}, /* 0x6c1a */
            {8'h00}, /* 0x6c19 */
            {8'h00}, /* 0x6c18 */
            {8'h00}, /* 0x6c17 */
            {8'h00}, /* 0x6c16 */
            {8'h00}, /* 0x6c15 */
            {8'h00}, /* 0x6c14 */
            {8'h00}, /* 0x6c13 */
            {8'h00}, /* 0x6c12 */
            {8'h00}, /* 0x6c11 */
            {8'h00}, /* 0x6c10 */
            {8'h00}, /* 0x6c0f */
            {8'h00}, /* 0x6c0e */
            {8'h00}, /* 0x6c0d */
            {8'h00}, /* 0x6c0c */
            {8'h00}, /* 0x6c0b */
            {8'h00}, /* 0x6c0a */
            {8'h00}, /* 0x6c09 */
            {8'h00}, /* 0x6c08 */
            {8'h00}, /* 0x6c07 */
            {8'h00}, /* 0x6c06 */
            {8'h00}, /* 0x6c05 */
            {8'h00}, /* 0x6c04 */
            {8'h00}, /* 0x6c03 */
            {8'h00}, /* 0x6c02 */
            {8'h00}, /* 0x6c01 */
            {8'h00}, /* 0x6c00 */
            {8'h00}, /* 0x6bff */
            {8'h00}, /* 0x6bfe */
            {8'h00}, /* 0x6bfd */
            {8'h00}, /* 0x6bfc */
            {8'h00}, /* 0x6bfb */
            {8'h00}, /* 0x6bfa */
            {8'h00}, /* 0x6bf9 */
            {8'h00}, /* 0x6bf8 */
            {8'h00}, /* 0x6bf7 */
            {8'h00}, /* 0x6bf6 */
            {8'h00}, /* 0x6bf5 */
            {8'h00}, /* 0x6bf4 */
            {8'h00}, /* 0x6bf3 */
            {8'h00}, /* 0x6bf2 */
            {8'h00}, /* 0x6bf1 */
            {8'h00}, /* 0x6bf0 */
            {8'h00}, /* 0x6bef */
            {8'h00}, /* 0x6bee */
            {8'h00}, /* 0x6bed */
            {8'h00}, /* 0x6bec */
            {8'h00}, /* 0x6beb */
            {8'h00}, /* 0x6bea */
            {8'h00}, /* 0x6be9 */
            {8'h00}, /* 0x6be8 */
            {8'h00}, /* 0x6be7 */
            {8'h00}, /* 0x6be6 */
            {8'h00}, /* 0x6be5 */
            {8'h00}, /* 0x6be4 */
            {8'h00}, /* 0x6be3 */
            {8'h00}, /* 0x6be2 */
            {8'h00}, /* 0x6be1 */
            {8'h00}, /* 0x6be0 */
            {8'h00}, /* 0x6bdf */
            {8'h00}, /* 0x6bde */
            {8'h00}, /* 0x6bdd */
            {8'h00}, /* 0x6bdc */
            {8'h00}, /* 0x6bdb */
            {8'h00}, /* 0x6bda */
            {8'h00}, /* 0x6bd9 */
            {8'h00}, /* 0x6bd8 */
            {8'h00}, /* 0x6bd7 */
            {8'h00}, /* 0x6bd6 */
            {8'h00}, /* 0x6bd5 */
            {8'h00}, /* 0x6bd4 */
            {8'h00}, /* 0x6bd3 */
            {8'h00}, /* 0x6bd2 */
            {8'h00}, /* 0x6bd1 */
            {8'h00}, /* 0x6bd0 */
            {8'h00}, /* 0x6bcf */
            {8'h00}, /* 0x6bce */
            {8'h00}, /* 0x6bcd */
            {8'h00}, /* 0x6bcc */
            {8'h00}, /* 0x6bcb */
            {8'h00}, /* 0x6bca */
            {8'h00}, /* 0x6bc9 */
            {8'h00}, /* 0x6bc8 */
            {8'h00}, /* 0x6bc7 */
            {8'h00}, /* 0x6bc6 */
            {8'h00}, /* 0x6bc5 */
            {8'h00}, /* 0x6bc4 */
            {8'h00}, /* 0x6bc3 */
            {8'h00}, /* 0x6bc2 */
            {8'h00}, /* 0x6bc1 */
            {8'h00}, /* 0x6bc0 */
            {8'h00}, /* 0x6bbf */
            {8'h00}, /* 0x6bbe */
            {8'h00}, /* 0x6bbd */
            {8'h00}, /* 0x6bbc */
            {8'h00}, /* 0x6bbb */
            {8'h00}, /* 0x6bba */
            {8'h00}, /* 0x6bb9 */
            {8'h00}, /* 0x6bb8 */
            {8'h00}, /* 0x6bb7 */
            {8'h00}, /* 0x6bb6 */
            {8'h00}, /* 0x6bb5 */
            {8'h00}, /* 0x6bb4 */
            {8'h00}, /* 0x6bb3 */
            {8'h00}, /* 0x6bb2 */
            {8'h00}, /* 0x6bb1 */
            {8'h00}, /* 0x6bb0 */
            {8'h00}, /* 0x6baf */
            {8'h00}, /* 0x6bae */
            {8'h00}, /* 0x6bad */
            {8'h00}, /* 0x6bac */
            {8'h00}, /* 0x6bab */
            {8'h00}, /* 0x6baa */
            {8'h00}, /* 0x6ba9 */
            {8'h00}, /* 0x6ba8 */
            {8'h00}, /* 0x6ba7 */
            {8'h00}, /* 0x6ba6 */
            {8'h00}, /* 0x6ba5 */
            {8'h00}, /* 0x6ba4 */
            {8'h00}, /* 0x6ba3 */
            {8'h00}, /* 0x6ba2 */
            {8'h00}, /* 0x6ba1 */
            {8'h00}, /* 0x6ba0 */
            {8'h00}, /* 0x6b9f */
            {8'h00}, /* 0x6b9e */
            {8'h00}, /* 0x6b9d */
            {8'h00}, /* 0x6b9c */
            {8'h00}, /* 0x6b9b */
            {8'h00}, /* 0x6b9a */
            {8'h00}, /* 0x6b99 */
            {8'h00}, /* 0x6b98 */
            {8'h00}, /* 0x6b97 */
            {8'h00}, /* 0x6b96 */
            {8'h00}, /* 0x6b95 */
            {8'h00}, /* 0x6b94 */
            {8'h00}, /* 0x6b93 */
            {8'h00}, /* 0x6b92 */
            {8'h00}, /* 0x6b91 */
            {8'h00}, /* 0x6b90 */
            {8'h00}, /* 0x6b8f */
            {8'h00}, /* 0x6b8e */
            {8'h00}, /* 0x6b8d */
            {8'h00}, /* 0x6b8c */
            {8'h00}, /* 0x6b8b */
            {8'h00}, /* 0x6b8a */
            {8'h00}, /* 0x6b89 */
            {8'h00}, /* 0x6b88 */
            {8'h00}, /* 0x6b87 */
            {8'h00}, /* 0x6b86 */
            {8'h00}, /* 0x6b85 */
            {8'h00}, /* 0x6b84 */
            {8'h00}, /* 0x6b83 */
            {8'h00}, /* 0x6b82 */
            {8'h00}, /* 0x6b81 */
            {8'h00}, /* 0x6b80 */
            {8'h00}, /* 0x6b7f */
            {8'h00}, /* 0x6b7e */
            {8'h00}, /* 0x6b7d */
            {8'h00}, /* 0x6b7c */
            {8'h00}, /* 0x6b7b */
            {8'h00}, /* 0x6b7a */
            {8'h00}, /* 0x6b79 */
            {8'h00}, /* 0x6b78 */
            {8'h00}, /* 0x6b77 */
            {8'h00}, /* 0x6b76 */
            {8'h00}, /* 0x6b75 */
            {8'h00}, /* 0x6b74 */
            {8'h00}, /* 0x6b73 */
            {8'h00}, /* 0x6b72 */
            {8'h00}, /* 0x6b71 */
            {8'h00}, /* 0x6b70 */
            {8'h00}, /* 0x6b6f */
            {8'h00}, /* 0x6b6e */
            {8'h00}, /* 0x6b6d */
            {8'h00}, /* 0x6b6c */
            {8'h00}, /* 0x6b6b */
            {8'h00}, /* 0x6b6a */
            {8'h00}, /* 0x6b69 */
            {8'h00}, /* 0x6b68 */
            {8'h00}, /* 0x6b67 */
            {8'h00}, /* 0x6b66 */
            {8'h00}, /* 0x6b65 */
            {8'h00}, /* 0x6b64 */
            {8'h00}, /* 0x6b63 */
            {8'h00}, /* 0x6b62 */
            {8'h00}, /* 0x6b61 */
            {8'h00}, /* 0x6b60 */
            {8'h00}, /* 0x6b5f */
            {8'h00}, /* 0x6b5e */
            {8'h00}, /* 0x6b5d */
            {8'h00}, /* 0x6b5c */
            {8'h00}, /* 0x6b5b */
            {8'h00}, /* 0x6b5a */
            {8'h00}, /* 0x6b59 */
            {8'h00}, /* 0x6b58 */
            {8'h00}, /* 0x6b57 */
            {8'h00}, /* 0x6b56 */
            {8'h00}, /* 0x6b55 */
            {8'h00}, /* 0x6b54 */
            {8'h00}, /* 0x6b53 */
            {8'h00}, /* 0x6b52 */
            {8'h00}, /* 0x6b51 */
            {8'h00}, /* 0x6b50 */
            {8'h00}, /* 0x6b4f */
            {8'h00}, /* 0x6b4e */
            {8'h00}, /* 0x6b4d */
            {8'h00}, /* 0x6b4c */
            {8'h00}, /* 0x6b4b */
            {8'h00}, /* 0x6b4a */
            {8'h00}, /* 0x6b49 */
            {8'h00}, /* 0x6b48 */
            {8'h00}, /* 0x6b47 */
            {8'h00}, /* 0x6b46 */
            {8'h00}, /* 0x6b45 */
            {8'h00}, /* 0x6b44 */
            {8'h00}, /* 0x6b43 */
            {8'h00}, /* 0x6b42 */
            {8'h00}, /* 0x6b41 */
            {8'h00}, /* 0x6b40 */
            {8'h00}, /* 0x6b3f */
            {8'h00}, /* 0x6b3e */
            {8'h00}, /* 0x6b3d */
            {8'h00}, /* 0x6b3c */
            {8'h00}, /* 0x6b3b */
            {8'h00}, /* 0x6b3a */
            {8'h00}, /* 0x6b39 */
            {8'h00}, /* 0x6b38 */
            {8'h00}, /* 0x6b37 */
            {8'h00}, /* 0x6b36 */
            {8'h00}, /* 0x6b35 */
            {8'h00}, /* 0x6b34 */
            {8'h00}, /* 0x6b33 */
            {8'h00}, /* 0x6b32 */
            {8'h00}, /* 0x6b31 */
            {8'h00}, /* 0x6b30 */
            {8'h00}, /* 0x6b2f */
            {8'h00}, /* 0x6b2e */
            {8'h00}, /* 0x6b2d */
            {8'h00}, /* 0x6b2c */
            {8'h00}, /* 0x6b2b */
            {8'h00}, /* 0x6b2a */
            {8'h00}, /* 0x6b29 */
            {8'h00}, /* 0x6b28 */
            {8'h00}, /* 0x6b27 */
            {8'h00}, /* 0x6b26 */
            {8'h00}, /* 0x6b25 */
            {8'h00}, /* 0x6b24 */
            {8'h00}, /* 0x6b23 */
            {8'h00}, /* 0x6b22 */
            {8'h00}, /* 0x6b21 */
            {8'h00}, /* 0x6b20 */
            {8'h00}, /* 0x6b1f */
            {8'h00}, /* 0x6b1e */
            {8'h00}, /* 0x6b1d */
            {8'h00}, /* 0x6b1c */
            {8'h00}, /* 0x6b1b */
            {8'h00}, /* 0x6b1a */
            {8'h00}, /* 0x6b19 */
            {8'h00}, /* 0x6b18 */
            {8'h00}, /* 0x6b17 */
            {8'h00}, /* 0x6b16 */
            {8'h00}, /* 0x6b15 */
            {8'h00}, /* 0x6b14 */
            {8'h00}, /* 0x6b13 */
            {8'h00}, /* 0x6b12 */
            {8'h00}, /* 0x6b11 */
            {8'h00}, /* 0x6b10 */
            {8'h00}, /* 0x6b0f */
            {8'h00}, /* 0x6b0e */
            {8'h00}, /* 0x6b0d */
            {8'h00}, /* 0x6b0c */
            {8'h00}, /* 0x6b0b */
            {8'h00}, /* 0x6b0a */
            {8'h00}, /* 0x6b09 */
            {8'h00}, /* 0x6b08 */
            {8'h00}, /* 0x6b07 */
            {8'h00}, /* 0x6b06 */
            {8'h00}, /* 0x6b05 */
            {8'h00}, /* 0x6b04 */
            {8'h00}, /* 0x6b03 */
            {8'h00}, /* 0x6b02 */
            {8'h00}, /* 0x6b01 */
            {8'h00}, /* 0x6b00 */
            {8'h00}, /* 0x6aff */
            {8'h00}, /* 0x6afe */
            {8'h00}, /* 0x6afd */
            {8'h00}, /* 0x6afc */
            {8'h00}, /* 0x6afb */
            {8'h00}, /* 0x6afa */
            {8'h00}, /* 0x6af9 */
            {8'h00}, /* 0x6af8 */
            {8'h00}, /* 0x6af7 */
            {8'h00}, /* 0x6af6 */
            {8'h00}, /* 0x6af5 */
            {8'h00}, /* 0x6af4 */
            {8'h00}, /* 0x6af3 */
            {8'h00}, /* 0x6af2 */
            {8'h00}, /* 0x6af1 */
            {8'h00}, /* 0x6af0 */
            {8'h00}, /* 0x6aef */
            {8'h00}, /* 0x6aee */
            {8'h00}, /* 0x6aed */
            {8'h00}, /* 0x6aec */
            {8'h00}, /* 0x6aeb */
            {8'h00}, /* 0x6aea */
            {8'h00}, /* 0x6ae9 */
            {8'h00}, /* 0x6ae8 */
            {8'h00}, /* 0x6ae7 */
            {8'h00}, /* 0x6ae6 */
            {8'h00}, /* 0x6ae5 */
            {8'h00}, /* 0x6ae4 */
            {8'h00}, /* 0x6ae3 */
            {8'h00}, /* 0x6ae2 */
            {8'h00}, /* 0x6ae1 */
            {8'h00}, /* 0x6ae0 */
            {8'h00}, /* 0x6adf */
            {8'h00}, /* 0x6ade */
            {8'h00}, /* 0x6add */
            {8'h00}, /* 0x6adc */
            {8'h00}, /* 0x6adb */
            {8'h00}, /* 0x6ada */
            {8'h00}, /* 0x6ad9 */
            {8'h00}, /* 0x6ad8 */
            {8'h00}, /* 0x6ad7 */
            {8'h00}, /* 0x6ad6 */
            {8'h00}, /* 0x6ad5 */
            {8'h00}, /* 0x6ad4 */
            {8'h00}, /* 0x6ad3 */
            {8'h00}, /* 0x6ad2 */
            {8'h00}, /* 0x6ad1 */
            {8'h00}, /* 0x6ad0 */
            {8'h00}, /* 0x6acf */
            {8'h00}, /* 0x6ace */
            {8'h00}, /* 0x6acd */
            {8'h00}, /* 0x6acc */
            {8'h00}, /* 0x6acb */
            {8'h00}, /* 0x6aca */
            {8'h00}, /* 0x6ac9 */
            {8'h00}, /* 0x6ac8 */
            {8'h00}, /* 0x6ac7 */
            {8'h00}, /* 0x6ac6 */
            {8'h00}, /* 0x6ac5 */
            {8'h00}, /* 0x6ac4 */
            {8'h00}, /* 0x6ac3 */
            {8'h00}, /* 0x6ac2 */
            {8'h00}, /* 0x6ac1 */
            {8'h00}, /* 0x6ac0 */
            {8'h00}, /* 0x6abf */
            {8'h00}, /* 0x6abe */
            {8'h00}, /* 0x6abd */
            {8'h00}, /* 0x6abc */
            {8'h00}, /* 0x6abb */
            {8'h00}, /* 0x6aba */
            {8'h00}, /* 0x6ab9 */
            {8'h00}, /* 0x6ab8 */
            {8'h00}, /* 0x6ab7 */
            {8'h00}, /* 0x6ab6 */
            {8'h00}, /* 0x6ab5 */
            {8'h00}, /* 0x6ab4 */
            {8'h00}, /* 0x6ab3 */
            {8'h00}, /* 0x6ab2 */
            {8'h00}, /* 0x6ab1 */
            {8'h00}, /* 0x6ab0 */
            {8'h00}, /* 0x6aaf */
            {8'h00}, /* 0x6aae */
            {8'h00}, /* 0x6aad */
            {8'h00}, /* 0x6aac */
            {8'h00}, /* 0x6aab */
            {8'h00}, /* 0x6aaa */
            {8'h00}, /* 0x6aa9 */
            {8'h00}, /* 0x6aa8 */
            {8'h00}, /* 0x6aa7 */
            {8'h00}, /* 0x6aa6 */
            {8'h00}, /* 0x6aa5 */
            {8'h00}, /* 0x6aa4 */
            {8'h00}, /* 0x6aa3 */
            {8'h00}, /* 0x6aa2 */
            {8'h00}, /* 0x6aa1 */
            {8'h00}, /* 0x6aa0 */
            {8'h00}, /* 0x6a9f */
            {8'h00}, /* 0x6a9e */
            {8'h00}, /* 0x6a9d */
            {8'h00}, /* 0x6a9c */
            {8'h00}, /* 0x6a9b */
            {8'h00}, /* 0x6a9a */
            {8'h00}, /* 0x6a99 */
            {8'h00}, /* 0x6a98 */
            {8'h00}, /* 0x6a97 */
            {8'h00}, /* 0x6a96 */
            {8'h00}, /* 0x6a95 */
            {8'h00}, /* 0x6a94 */
            {8'h00}, /* 0x6a93 */
            {8'h00}, /* 0x6a92 */
            {8'h00}, /* 0x6a91 */
            {8'h00}, /* 0x6a90 */
            {8'h00}, /* 0x6a8f */
            {8'h00}, /* 0x6a8e */
            {8'h00}, /* 0x6a8d */
            {8'h00}, /* 0x6a8c */
            {8'h00}, /* 0x6a8b */
            {8'h00}, /* 0x6a8a */
            {8'h00}, /* 0x6a89 */
            {8'h00}, /* 0x6a88 */
            {8'h00}, /* 0x6a87 */
            {8'h00}, /* 0x6a86 */
            {8'h00}, /* 0x6a85 */
            {8'h00}, /* 0x6a84 */
            {8'h00}, /* 0x6a83 */
            {8'h00}, /* 0x6a82 */
            {8'h00}, /* 0x6a81 */
            {8'h00}, /* 0x6a80 */
            {8'h00}, /* 0x6a7f */
            {8'h00}, /* 0x6a7e */
            {8'h00}, /* 0x6a7d */
            {8'h00}, /* 0x6a7c */
            {8'h00}, /* 0x6a7b */
            {8'h00}, /* 0x6a7a */
            {8'h00}, /* 0x6a79 */
            {8'h00}, /* 0x6a78 */
            {8'h00}, /* 0x6a77 */
            {8'h00}, /* 0x6a76 */
            {8'h00}, /* 0x6a75 */
            {8'h00}, /* 0x6a74 */
            {8'h00}, /* 0x6a73 */
            {8'h00}, /* 0x6a72 */
            {8'h00}, /* 0x6a71 */
            {8'h00}, /* 0x6a70 */
            {8'h00}, /* 0x6a6f */
            {8'h00}, /* 0x6a6e */
            {8'h00}, /* 0x6a6d */
            {8'h00}, /* 0x6a6c */
            {8'h00}, /* 0x6a6b */
            {8'h00}, /* 0x6a6a */
            {8'h00}, /* 0x6a69 */
            {8'h00}, /* 0x6a68 */
            {8'h00}, /* 0x6a67 */
            {8'h00}, /* 0x6a66 */
            {8'h00}, /* 0x6a65 */
            {8'h00}, /* 0x6a64 */
            {8'h00}, /* 0x6a63 */
            {8'h00}, /* 0x6a62 */
            {8'h00}, /* 0x6a61 */
            {8'h00}, /* 0x6a60 */
            {8'h00}, /* 0x6a5f */
            {8'h00}, /* 0x6a5e */
            {8'h00}, /* 0x6a5d */
            {8'h00}, /* 0x6a5c */
            {8'h00}, /* 0x6a5b */
            {8'h00}, /* 0x6a5a */
            {8'h00}, /* 0x6a59 */
            {8'h00}, /* 0x6a58 */
            {8'h00}, /* 0x6a57 */
            {8'h00}, /* 0x6a56 */
            {8'h00}, /* 0x6a55 */
            {8'h00}, /* 0x6a54 */
            {8'h00}, /* 0x6a53 */
            {8'h00}, /* 0x6a52 */
            {8'h00}, /* 0x6a51 */
            {8'h00}, /* 0x6a50 */
            {8'h00}, /* 0x6a4f */
            {8'h00}, /* 0x6a4e */
            {8'h00}, /* 0x6a4d */
            {8'h00}, /* 0x6a4c */
            {8'h00}, /* 0x6a4b */
            {8'h00}, /* 0x6a4a */
            {8'h00}, /* 0x6a49 */
            {8'h00}, /* 0x6a48 */
            {8'h00}, /* 0x6a47 */
            {8'h00}, /* 0x6a46 */
            {8'h00}, /* 0x6a45 */
            {8'h00}, /* 0x6a44 */
            {8'h00}, /* 0x6a43 */
            {8'h00}, /* 0x6a42 */
            {8'h00}, /* 0x6a41 */
            {8'h00}, /* 0x6a40 */
            {8'h00}, /* 0x6a3f */
            {8'h00}, /* 0x6a3e */
            {8'h00}, /* 0x6a3d */
            {8'h00}, /* 0x6a3c */
            {8'h00}, /* 0x6a3b */
            {8'h00}, /* 0x6a3a */
            {8'h00}, /* 0x6a39 */
            {8'h00}, /* 0x6a38 */
            {8'h00}, /* 0x6a37 */
            {8'h00}, /* 0x6a36 */
            {8'h00}, /* 0x6a35 */
            {8'h00}, /* 0x6a34 */
            {8'h00}, /* 0x6a33 */
            {8'h00}, /* 0x6a32 */
            {8'h00}, /* 0x6a31 */
            {8'h00}, /* 0x6a30 */
            {8'h00}, /* 0x6a2f */
            {8'h00}, /* 0x6a2e */
            {8'h00}, /* 0x6a2d */
            {8'h00}, /* 0x6a2c */
            {8'h00}, /* 0x6a2b */
            {8'h00}, /* 0x6a2a */
            {8'h00}, /* 0x6a29 */
            {8'h00}, /* 0x6a28 */
            {8'h00}, /* 0x6a27 */
            {8'h00}, /* 0x6a26 */
            {8'h00}, /* 0x6a25 */
            {8'h00}, /* 0x6a24 */
            {8'h00}, /* 0x6a23 */
            {8'h00}, /* 0x6a22 */
            {8'h00}, /* 0x6a21 */
            {8'h00}, /* 0x6a20 */
            {8'h00}, /* 0x6a1f */
            {8'h00}, /* 0x6a1e */
            {8'h00}, /* 0x6a1d */
            {8'h00}, /* 0x6a1c */
            {8'h00}, /* 0x6a1b */
            {8'h00}, /* 0x6a1a */
            {8'h00}, /* 0x6a19 */
            {8'h00}, /* 0x6a18 */
            {8'h00}, /* 0x6a17 */
            {8'h00}, /* 0x6a16 */
            {8'h00}, /* 0x6a15 */
            {8'h00}, /* 0x6a14 */
            {8'h00}, /* 0x6a13 */
            {8'h00}, /* 0x6a12 */
            {8'h00}, /* 0x6a11 */
            {8'h00}, /* 0x6a10 */
            {8'h00}, /* 0x6a0f */
            {8'h00}, /* 0x6a0e */
            {8'h00}, /* 0x6a0d */
            {8'h00}, /* 0x6a0c */
            {8'h00}, /* 0x6a0b */
            {8'h00}, /* 0x6a0a */
            {8'h00}, /* 0x6a09 */
            {8'h00}, /* 0x6a08 */
            {8'h00}, /* 0x6a07 */
            {8'h00}, /* 0x6a06 */
            {8'h00}, /* 0x6a05 */
            {8'h00}, /* 0x6a04 */
            {8'h00}, /* 0x6a03 */
            {8'h00}, /* 0x6a02 */
            {8'h00}, /* 0x6a01 */
            {8'h00}, /* 0x6a00 */
            {8'h00}, /* 0x69ff */
            {8'h00}, /* 0x69fe */
            {8'h00}, /* 0x69fd */
            {8'h00}, /* 0x69fc */
            {8'h00}, /* 0x69fb */
            {8'h00}, /* 0x69fa */
            {8'h00}, /* 0x69f9 */
            {8'h00}, /* 0x69f8 */
            {8'h00}, /* 0x69f7 */
            {8'h00}, /* 0x69f6 */
            {8'h00}, /* 0x69f5 */
            {8'h00}, /* 0x69f4 */
            {8'h00}, /* 0x69f3 */
            {8'h00}, /* 0x69f2 */
            {8'h00}, /* 0x69f1 */
            {8'h00}, /* 0x69f0 */
            {8'h00}, /* 0x69ef */
            {8'h00}, /* 0x69ee */
            {8'h00}, /* 0x69ed */
            {8'h00}, /* 0x69ec */
            {8'h00}, /* 0x69eb */
            {8'h00}, /* 0x69ea */
            {8'h00}, /* 0x69e9 */
            {8'h00}, /* 0x69e8 */
            {8'h00}, /* 0x69e7 */
            {8'h00}, /* 0x69e6 */
            {8'h00}, /* 0x69e5 */
            {8'h00}, /* 0x69e4 */
            {8'h00}, /* 0x69e3 */
            {8'h00}, /* 0x69e2 */
            {8'h00}, /* 0x69e1 */
            {8'h00}, /* 0x69e0 */
            {8'h00}, /* 0x69df */
            {8'h00}, /* 0x69de */
            {8'h00}, /* 0x69dd */
            {8'h00}, /* 0x69dc */
            {8'h00}, /* 0x69db */
            {8'h00}, /* 0x69da */
            {8'h00}, /* 0x69d9 */
            {8'h00}, /* 0x69d8 */
            {8'h00}, /* 0x69d7 */
            {8'h00}, /* 0x69d6 */
            {8'h00}, /* 0x69d5 */
            {8'h00}, /* 0x69d4 */
            {8'h00}, /* 0x69d3 */
            {8'h00}, /* 0x69d2 */
            {8'h00}, /* 0x69d1 */
            {8'h00}, /* 0x69d0 */
            {8'h00}, /* 0x69cf */
            {8'h00}, /* 0x69ce */
            {8'h00}, /* 0x69cd */
            {8'h00}, /* 0x69cc */
            {8'h00}, /* 0x69cb */
            {8'h00}, /* 0x69ca */
            {8'h00}, /* 0x69c9 */
            {8'h00}, /* 0x69c8 */
            {8'h00}, /* 0x69c7 */
            {8'h00}, /* 0x69c6 */
            {8'h00}, /* 0x69c5 */
            {8'h00}, /* 0x69c4 */
            {8'h00}, /* 0x69c3 */
            {8'h00}, /* 0x69c2 */
            {8'h00}, /* 0x69c1 */
            {8'h00}, /* 0x69c0 */
            {8'h00}, /* 0x69bf */
            {8'h00}, /* 0x69be */
            {8'h00}, /* 0x69bd */
            {8'h00}, /* 0x69bc */
            {8'h00}, /* 0x69bb */
            {8'h00}, /* 0x69ba */
            {8'h00}, /* 0x69b9 */
            {8'h00}, /* 0x69b8 */
            {8'h00}, /* 0x69b7 */
            {8'h00}, /* 0x69b6 */
            {8'h00}, /* 0x69b5 */
            {8'h00}, /* 0x69b4 */
            {8'h00}, /* 0x69b3 */
            {8'h00}, /* 0x69b2 */
            {8'h00}, /* 0x69b1 */
            {8'h00}, /* 0x69b0 */
            {8'h00}, /* 0x69af */
            {8'h00}, /* 0x69ae */
            {8'h00}, /* 0x69ad */
            {8'h00}, /* 0x69ac */
            {8'h00}, /* 0x69ab */
            {8'h00}, /* 0x69aa */
            {8'h00}, /* 0x69a9 */
            {8'h00}, /* 0x69a8 */
            {8'h00}, /* 0x69a7 */
            {8'h00}, /* 0x69a6 */
            {8'h00}, /* 0x69a5 */
            {8'h00}, /* 0x69a4 */
            {8'h00}, /* 0x69a3 */
            {8'h00}, /* 0x69a2 */
            {8'h00}, /* 0x69a1 */
            {8'h00}, /* 0x69a0 */
            {8'h00}, /* 0x699f */
            {8'h00}, /* 0x699e */
            {8'h00}, /* 0x699d */
            {8'h00}, /* 0x699c */
            {8'h00}, /* 0x699b */
            {8'h00}, /* 0x699a */
            {8'h00}, /* 0x6999 */
            {8'h00}, /* 0x6998 */
            {8'h00}, /* 0x6997 */
            {8'h00}, /* 0x6996 */
            {8'h00}, /* 0x6995 */
            {8'h00}, /* 0x6994 */
            {8'h00}, /* 0x6993 */
            {8'h00}, /* 0x6992 */
            {8'h00}, /* 0x6991 */
            {8'h00}, /* 0x6990 */
            {8'h00}, /* 0x698f */
            {8'h00}, /* 0x698e */
            {8'h00}, /* 0x698d */
            {8'h00}, /* 0x698c */
            {8'h00}, /* 0x698b */
            {8'h00}, /* 0x698a */
            {8'h00}, /* 0x6989 */
            {8'h00}, /* 0x6988 */
            {8'h00}, /* 0x6987 */
            {8'h00}, /* 0x6986 */
            {8'h00}, /* 0x6985 */
            {8'h00}, /* 0x6984 */
            {8'h00}, /* 0x6983 */
            {8'h00}, /* 0x6982 */
            {8'h00}, /* 0x6981 */
            {8'h00}, /* 0x6980 */
            {8'h00}, /* 0x697f */
            {8'h00}, /* 0x697e */
            {8'h00}, /* 0x697d */
            {8'h00}, /* 0x697c */
            {8'h00}, /* 0x697b */
            {8'h00}, /* 0x697a */
            {8'h00}, /* 0x6979 */
            {8'h00}, /* 0x6978 */
            {8'h00}, /* 0x6977 */
            {8'h00}, /* 0x6976 */
            {8'h00}, /* 0x6975 */
            {8'h00}, /* 0x6974 */
            {8'h00}, /* 0x6973 */
            {8'h00}, /* 0x6972 */
            {8'h00}, /* 0x6971 */
            {8'h00}, /* 0x6970 */
            {8'h00}, /* 0x696f */
            {8'h00}, /* 0x696e */
            {8'h00}, /* 0x696d */
            {8'h00}, /* 0x696c */
            {8'h00}, /* 0x696b */
            {8'h00}, /* 0x696a */
            {8'h00}, /* 0x6969 */
            {8'h00}, /* 0x6968 */
            {8'h00}, /* 0x6967 */
            {8'h00}, /* 0x6966 */
            {8'h00}, /* 0x6965 */
            {8'h00}, /* 0x6964 */
            {8'h00}, /* 0x6963 */
            {8'h00}, /* 0x6962 */
            {8'h00}, /* 0x6961 */
            {8'h00}, /* 0x6960 */
            {8'h00}, /* 0x695f */
            {8'h00}, /* 0x695e */
            {8'h00}, /* 0x695d */
            {8'h00}, /* 0x695c */
            {8'h00}, /* 0x695b */
            {8'h00}, /* 0x695a */
            {8'h00}, /* 0x6959 */
            {8'h00}, /* 0x6958 */
            {8'h00}, /* 0x6957 */
            {8'h00}, /* 0x6956 */
            {8'h00}, /* 0x6955 */
            {8'h00}, /* 0x6954 */
            {8'h00}, /* 0x6953 */
            {8'h00}, /* 0x6952 */
            {8'h00}, /* 0x6951 */
            {8'h00}, /* 0x6950 */
            {8'h00}, /* 0x694f */
            {8'h00}, /* 0x694e */
            {8'h00}, /* 0x694d */
            {8'h00}, /* 0x694c */
            {8'h00}, /* 0x694b */
            {8'h00}, /* 0x694a */
            {8'h00}, /* 0x6949 */
            {8'h00}, /* 0x6948 */
            {8'h00}, /* 0x6947 */
            {8'h00}, /* 0x6946 */
            {8'h00}, /* 0x6945 */
            {8'h00}, /* 0x6944 */
            {8'h00}, /* 0x6943 */
            {8'h00}, /* 0x6942 */
            {8'h00}, /* 0x6941 */
            {8'h00}, /* 0x6940 */
            {8'h00}, /* 0x693f */
            {8'h00}, /* 0x693e */
            {8'h00}, /* 0x693d */
            {8'h00}, /* 0x693c */
            {8'h00}, /* 0x693b */
            {8'h00}, /* 0x693a */
            {8'h00}, /* 0x6939 */
            {8'h00}, /* 0x6938 */
            {8'h00}, /* 0x6937 */
            {8'h00}, /* 0x6936 */
            {8'h00}, /* 0x6935 */
            {8'h00}, /* 0x6934 */
            {8'h00}, /* 0x6933 */
            {8'h00}, /* 0x6932 */
            {8'h00}, /* 0x6931 */
            {8'h00}, /* 0x6930 */
            {8'h00}, /* 0x692f */
            {8'h00}, /* 0x692e */
            {8'h00}, /* 0x692d */
            {8'h00}, /* 0x692c */
            {8'h00}, /* 0x692b */
            {8'h00}, /* 0x692a */
            {8'h00}, /* 0x6929 */
            {8'h00}, /* 0x6928 */
            {8'h00}, /* 0x6927 */
            {8'h00}, /* 0x6926 */
            {8'h00}, /* 0x6925 */
            {8'h00}, /* 0x6924 */
            {8'h00}, /* 0x6923 */
            {8'h00}, /* 0x6922 */
            {8'h00}, /* 0x6921 */
            {8'h00}, /* 0x6920 */
            {8'h00}, /* 0x691f */
            {8'h00}, /* 0x691e */
            {8'h00}, /* 0x691d */
            {8'h00}, /* 0x691c */
            {8'h00}, /* 0x691b */
            {8'h00}, /* 0x691a */
            {8'h00}, /* 0x6919 */
            {8'h00}, /* 0x6918 */
            {8'h00}, /* 0x6917 */
            {8'h00}, /* 0x6916 */
            {8'h00}, /* 0x6915 */
            {8'h00}, /* 0x6914 */
            {8'h00}, /* 0x6913 */
            {8'h00}, /* 0x6912 */
            {8'h00}, /* 0x6911 */
            {8'h00}, /* 0x6910 */
            {8'h00}, /* 0x690f */
            {8'h00}, /* 0x690e */
            {8'h00}, /* 0x690d */
            {8'h00}, /* 0x690c */
            {8'h00}, /* 0x690b */
            {8'h00}, /* 0x690a */
            {8'h00}, /* 0x6909 */
            {8'h00}, /* 0x6908 */
            {8'h00}, /* 0x6907 */
            {8'h00}, /* 0x6906 */
            {8'h00}, /* 0x6905 */
            {8'h00}, /* 0x6904 */
            {8'h00}, /* 0x6903 */
            {8'h00}, /* 0x6902 */
            {8'h00}, /* 0x6901 */
            {8'h00}, /* 0x6900 */
            {8'h00}, /* 0x68ff */
            {8'h00}, /* 0x68fe */
            {8'h00}, /* 0x68fd */
            {8'h00}, /* 0x68fc */
            {8'h00}, /* 0x68fb */
            {8'h00}, /* 0x68fa */
            {8'h00}, /* 0x68f9 */
            {8'h00}, /* 0x68f8 */
            {8'h00}, /* 0x68f7 */
            {8'h00}, /* 0x68f6 */
            {8'h00}, /* 0x68f5 */
            {8'h00}, /* 0x68f4 */
            {8'h00}, /* 0x68f3 */
            {8'h00}, /* 0x68f2 */
            {8'h00}, /* 0x68f1 */
            {8'h00}, /* 0x68f0 */
            {8'h00}, /* 0x68ef */
            {8'h00}, /* 0x68ee */
            {8'h00}, /* 0x68ed */
            {8'h00}, /* 0x68ec */
            {8'h00}, /* 0x68eb */
            {8'h00}, /* 0x68ea */
            {8'h00}, /* 0x68e9 */
            {8'h00}, /* 0x68e8 */
            {8'h00}, /* 0x68e7 */
            {8'h00}, /* 0x68e6 */
            {8'h00}, /* 0x68e5 */
            {8'h00}, /* 0x68e4 */
            {8'h00}, /* 0x68e3 */
            {8'h00}, /* 0x68e2 */
            {8'h00}, /* 0x68e1 */
            {8'h00}, /* 0x68e0 */
            {8'h00}, /* 0x68df */
            {8'h00}, /* 0x68de */
            {8'h00}, /* 0x68dd */
            {8'h00}, /* 0x68dc */
            {8'h00}, /* 0x68db */
            {8'h00}, /* 0x68da */
            {8'h00}, /* 0x68d9 */
            {8'h00}, /* 0x68d8 */
            {8'h00}, /* 0x68d7 */
            {8'h00}, /* 0x68d6 */
            {8'h00}, /* 0x68d5 */
            {8'h00}, /* 0x68d4 */
            {8'h00}, /* 0x68d3 */
            {8'h00}, /* 0x68d2 */
            {8'h00}, /* 0x68d1 */
            {8'h00}, /* 0x68d0 */
            {8'h00}, /* 0x68cf */
            {8'h00}, /* 0x68ce */
            {8'h00}, /* 0x68cd */
            {8'h00}, /* 0x68cc */
            {8'h00}, /* 0x68cb */
            {8'h00}, /* 0x68ca */
            {8'h00}, /* 0x68c9 */
            {8'h00}, /* 0x68c8 */
            {8'h00}, /* 0x68c7 */
            {8'h00}, /* 0x68c6 */
            {8'h00}, /* 0x68c5 */
            {8'h00}, /* 0x68c4 */
            {8'h00}, /* 0x68c3 */
            {8'h00}, /* 0x68c2 */
            {8'h00}, /* 0x68c1 */
            {8'h00}, /* 0x68c0 */
            {8'h00}, /* 0x68bf */
            {8'h00}, /* 0x68be */
            {8'h00}, /* 0x68bd */
            {8'h00}, /* 0x68bc */
            {8'h00}, /* 0x68bb */
            {8'h00}, /* 0x68ba */
            {8'h00}, /* 0x68b9 */
            {8'h00}, /* 0x68b8 */
            {8'h00}, /* 0x68b7 */
            {8'h00}, /* 0x68b6 */
            {8'h00}, /* 0x68b5 */
            {8'h00}, /* 0x68b4 */
            {8'h00}, /* 0x68b3 */
            {8'h00}, /* 0x68b2 */
            {8'h00}, /* 0x68b1 */
            {8'h00}, /* 0x68b0 */
            {8'h00}, /* 0x68af */
            {8'h00}, /* 0x68ae */
            {8'h00}, /* 0x68ad */
            {8'h00}, /* 0x68ac */
            {8'h00}, /* 0x68ab */
            {8'h00}, /* 0x68aa */
            {8'h00}, /* 0x68a9 */
            {8'h00}, /* 0x68a8 */
            {8'h00}, /* 0x68a7 */
            {8'h00}, /* 0x68a6 */
            {8'h00}, /* 0x68a5 */
            {8'h00}, /* 0x68a4 */
            {8'h00}, /* 0x68a3 */
            {8'h00}, /* 0x68a2 */
            {8'h00}, /* 0x68a1 */
            {8'h00}, /* 0x68a0 */
            {8'h00}, /* 0x689f */
            {8'h00}, /* 0x689e */
            {8'h00}, /* 0x689d */
            {8'h00}, /* 0x689c */
            {8'h00}, /* 0x689b */
            {8'h00}, /* 0x689a */
            {8'h00}, /* 0x6899 */
            {8'h00}, /* 0x6898 */
            {8'h00}, /* 0x6897 */
            {8'h00}, /* 0x6896 */
            {8'h00}, /* 0x6895 */
            {8'h00}, /* 0x6894 */
            {8'h00}, /* 0x6893 */
            {8'h00}, /* 0x6892 */
            {8'h00}, /* 0x6891 */
            {8'h00}, /* 0x6890 */
            {8'h00}, /* 0x688f */
            {8'h00}, /* 0x688e */
            {8'h00}, /* 0x688d */
            {8'h00}, /* 0x688c */
            {8'h00}, /* 0x688b */
            {8'h00}, /* 0x688a */
            {8'h00}, /* 0x6889 */
            {8'h00}, /* 0x6888 */
            {8'h00}, /* 0x6887 */
            {8'h00}, /* 0x6886 */
            {8'h00}, /* 0x6885 */
            {8'h00}, /* 0x6884 */
            {8'h00}, /* 0x6883 */
            {8'h00}, /* 0x6882 */
            {8'h00}, /* 0x6881 */
            {8'h00}, /* 0x6880 */
            {8'h00}, /* 0x687f */
            {8'h00}, /* 0x687e */
            {8'h00}, /* 0x687d */
            {8'h00}, /* 0x687c */
            {8'h00}, /* 0x687b */
            {8'h00}, /* 0x687a */
            {8'h00}, /* 0x6879 */
            {8'h00}, /* 0x6878 */
            {8'h00}, /* 0x6877 */
            {8'h00}, /* 0x6876 */
            {8'h00}, /* 0x6875 */
            {8'h00}, /* 0x6874 */
            {8'h00}, /* 0x6873 */
            {8'h00}, /* 0x6872 */
            {8'h00}, /* 0x6871 */
            {8'h00}, /* 0x6870 */
            {8'h00}, /* 0x686f */
            {8'h00}, /* 0x686e */
            {8'h00}, /* 0x686d */
            {8'h00}, /* 0x686c */
            {8'h00}, /* 0x686b */
            {8'h00}, /* 0x686a */
            {8'h00}, /* 0x6869 */
            {8'h00}, /* 0x6868 */
            {8'h00}, /* 0x6867 */
            {8'h00}, /* 0x6866 */
            {8'h00}, /* 0x6865 */
            {8'h00}, /* 0x6864 */
            {8'h00}, /* 0x6863 */
            {8'h00}, /* 0x6862 */
            {8'h00}, /* 0x6861 */
            {8'h00}, /* 0x6860 */
            {8'h00}, /* 0x685f */
            {8'h00}, /* 0x685e */
            {8'h00}, /* 0x685d */
            {8'h00}, /* 0x685c */
            {8'h00}, /* 0x685b */
            {8'h00}, /* 0x685a */
            {8'h00}, /* 0x6859 */
            {8'h00}, /* 0x6858 */
            {8'h00}, /* 0x6857 */
            {8'h00}, /* 0x6856 */
            {8'h00}, /* 0x6855 */
            {8'h00}, /* 0x6854 */
            {8'h00}, /* 0x6853 */
            {8'h00}, /* 0x6852 */
            {8'h00}, /* 0x6851 */
            {8'h00}, /* 0x6850 */
            {8'h00}, /* 0x684f */
            {8'h00}, /* 0x684e */
            {8'h00}, /* 0x684d */
            {8'h00}, /* 0x684c */
            {8'h00}, /* 0x684b */
            {8'h00}, /* 0x684a */
            {8'h00}, /* 0x6849 */
            {8'h00}, /* 0x6848 */
            {8'h00}, /* 0x6847 */
            {8'h00}, /* 0x6846 */
            {8'h00}, /* 0x6845 */
            {8'h00}, /* 0x6844 */
            {8'h00}, /* 0x6843 */
            {8'h00}, /* 0x6842 */
            {8'h00}, /* 0x6841 */
            {8'h00}, /* 0x6840 */
            {8'h00}, /* 0x683f */
            {8'h00}, /* 0x683e */
            {8'h00}, /* 0x683d */
            {8'h00}, /* 0x683c */
            {8'h00}, /* 0x683b */
            {8'h00}, /* 0x683a */
            {8'h00}, /* 0x6839 */
            {8'h00}, /* 0x6838 */
            {8'h00}, /* 0x6837 */
            {8'h00}, /* 0x6836 */
            {8'h00}, /* 0x6835 */
            {8'h00}, /* 0x6834 */
            {8'h00}, /* 0x6833 */
            {8'h00}, /* 0x6832 */
            {8'h00}, /* 0x6831 */
            {8'h00}, /* 0x6830 */
            {8'h00}, /* 0x682f */
            {8'h00}, /* 0x682e */
            {8'h00}, /* 0x682d */
            {8'h00}, /* 0x682c */
            {8'h00}, /* 0x682b */
            {8'h00}, /* 0x682a */
            {8'h00}, /* 0x6829 */
            {8'h00}, /* 0x6828 */
            {8'h00}, /* 0x6827 */
            {8'h00}, /* 0x6826 */
            {8'h00}, /* 0x6825 */
            {8'h00}, /* 0x6824 */
            {8'h00}, /* 0x6823 */
            {8'h00}, /* 0x6822 */
            {8'h00}, /* 0x6821 */
            {8'h00}, /* 0x6820 */
            {8'h00}, /* 0x681f */
            {8'h00}, /* 0x681e */
            {8'h00}, /* 0x681d */
            {8'h00}, /* 0x681c */
            {8'h00}, /* 0x681b */
            {8'h00}, /* 0x681a */
            {8'h00}, /* 0x6819 */
            {8'h00}, /* 0x6818 */
            {8'h00}, /* 0x6817 */
            {8'h00}, /* 0x6816 */
            {8'h00}, /* 0x6815 */
            {8'h00}, /* 0x6814 */
            {8'h00}, /* 0x6813 */
            {8'h00}, /* 0x6812 */
            {8'h00}, /* 0x6811 */
            {8'h00}, /* 0x6810 */
            {8'h00}, /* 0x680f */
            {8'h00}, /* 0x680e */
            {8'h00}, /* 0x680d */
            {8'h00}, /* 0x680c */
            {8'h00}, /* 0x680b */
            {8'h00}, /* 0x680a */
            {8'h00}, /* 0x6809 */
            {8'h00}, /* 0x6808 */
            {8'h00}, /* 0x6807 */
            {8'h00}, /* 0x6806 */
            {8'h00}, /* 0x6805 */
            {8'h00}, /* 0x6804 */
            {8'h00}, /* 0x6803 */
            {8'h00}, /* 0x6802 */
            {8'h00}, /* 0x6801 */
            {8'h00}, /* 0x6800 */
            {8'h00}, /* 0x67ff */
            {8'h00}, /* 0x67fe */
            {8'h00}, /* 0x67fd */
            {8'h00}, /* 0x67fc */
            {8'h00}, /* 0x67fb */
            {8'h00}, /* 0x67fa */
            {8'h00}, /* 0x67f9 */
            {8'h00}, /* 0x67f8 */
            {8'h00}, /* 0x67f7 */
            {8'h00}, /* 0x67f6 */
            {8'h00}, /* 0x67f5 */
            {8'h00}, /* 0x67f4 */
            {8'h00}, /* 0x67f3 */
            {8'h00}, /* 0x67f2 */
            {8'h00}, /* 0x67f1 */
            {8'h00}, /* 0x67f0 */
            {8'h00}, /* 0x67ef */
            {8'h00}, /* 0x67ee */
            {8'h00}, /* 0x67ed */
            {8'h00}, /* 0x67ec */
            {8'h00}, /* 0x67eb */
            {8'h00}, /* 0x67ea */
            {8'h00}, /* 0x67e9 */
            {8'h00}, /* 0x67e8 */
            {8'h00}, /* 0x67e7 */
            {8'h00}, /* 0x67e6 */
            {8'h00}, /* 0x67e5 */
            {8'h00}, /* 0x67e4 */
            {8'h00}, /* 0x67e3 */
            {8'h00}, /* 0x67e2 */
            {8'h00}, /* 0x67e1 */
            {8'h00}, /* 0x67e0 */
            {8'h00}, /* 0x67df */
            {8'h00}, /* 0x67de */
            {8'h00}, /* 0x67dd */
            {8'h00}, /* 0x67dc */
            {8'h00}, /* 0x67db */
            {8'h00}, /* 0x67da */
            {8'h00}, /* 0x67d9 */
            {8'h00}, /* 0x67d8 */
            {8'h00}, /* 0x67d7 */
            {8'h00}, /* 0x67d6 */
            {8'h00}, /* 0x67d5 */
            {8'h00}, /* 0x67d4 */
            {8'h00}, /* 0x67d3 */
            {8'h00}, /* 0x67d2 */
            {8'h00}, /* 0x67d1 */
            {8'h00}, /* 0x67d0 */
            {8'h00}, /* 0x67cf */
            {8'h00}, /* 0x67ce */
            {8'h00}, /* 0x67cd */
            {8'h00}, /* 0x67cc */
            {8'h00}, /* 0x67cb */
            {8'h00}, /* 0x67ca */
            {8'h00}, /* 0x67c9 */
            {8'h00}, /* 0x67c8 */
            {8'h00}, /* 0x67c7 */
            {8'h00}, /* 0x67c6 */
            {8'h00}, /* 0x67c5 */
            {8'h00}, /* 0x67c4 */
            {8'h00}, /* 0x67c3 */
            {8'h00}, /* 0x67c2 */
            {8'h00}, /* 0x67c1 */
            {8'h00}, /* 0x67c0 */
            {8'h00}, /* 0x67bf */
            {8'h00}, /* 0x67be */
            {8'h00}, /* 0x67bd */
            {8'h00}, /* 0x67bc */
            {8'h00}, /* 0x67bb */
            {8'h00}, /* 0x67ba */
            {8'h00}, /* 0x67b9 */
            {8'h00}, /* 0x67b8 */
            {8'h00}, /* 0x67b7 */
            {8'h00}, /* 0x67b6 */
            {8'h00}, /* 0x67b5 */
            {8'h00}, /* 0x67b4 */
            {8'h00}, /* 0x67b3 */
            {8'h00}, /* 0x67b2 */
            {8'h00}, /* 0x67b1 */
            {8'h00}, /* 0x67b0 */
            {8'h00}, /* 0x67af */
            {8'h00}, /* 0x67ae */
            {8'h00}, /* 0x67ad */
            {8'h00}, /* 0x67ac */
            {8'h00}, /* 0x67ab */
            {8'h00}, /* 0x67aa */
            {8'h00}, /* 0x67a9 */
            {8'h00}, /* 0x67a8 */
            {8'h00}, /* 0x67a7 */
            {8'h00}, /* 0x67a6 */
            {8'h00}, /* 0x67a5 */
            {8'h00}, /* 0x67a4 */
            {8'h00}, /* 0x67a3 */
            {8'h00}, /* 0x67a2 */
            {8'h00}, /* 0x67a1 */
            {8'h00}, /* 0x67a0 */
            {8'h00}, /* 0x679f */
            {8'h00}, /* 0x679e */
            {8'h00}, /* 0x679d */
            {8'h00}, /* 0x679c */
            {8'h00}, /* 0x679b */
            {8'h00}, /* 0x679a */
            {8'h00}, /* 0x6799 */
            {8'h00}, /* 0x6798 */
            {8'h00}, /* 0x6797 */
            {8'h00}, /* 0x6796 */
            {8'h00}, /* 0x6795 */
            {8'h00}, /* 0x6794 */
            {8'h00}, /* 0x6793 */
            {8'h00}, /* 0x6792 */
            {8'h00}, /* 0x6791 */
            {8'h00}, /* 0x6790 */
            {8'h00}, /* 0x678f */
            {8'h00}, /* 0x678e */
            {8'h00}, /* 0x678d */
            {8'h00}, /* 0x678c */
            {8'h00}, /* 0x678b */
            {8'h00}, /* 0x678a */
            {8'h00}, /* 0x6789 */
            {8'h00}, /* 0x6788 */
            {8'h00}, /* 0x6787 */
            {8'h00}, /* 0x6786 */
            {8'h00}, /* 0x6785 */
            {8'h00}, /* 0x6784 */
            {8'h00}, /* 0x6783 */
            {8'h00}, /* 0x6782 */
            {8'h00}, /* 0x6781 */
            {8'h00}, /* 0x6780 */
            {8'h00}, /* 0x677f */
            {8'h00}, /* 0x677e */
            {8'h00}, /* 0x677d */
            {8'h00}, /* 0x677c */
            {8'h00}, /* 0x677b */
            {8'h00}, /* 0x677a */
            {8'h00}, /* 0x6779 */
            {8'h00}, /* 0x6778 */
            {8'h00}, /* 0x6777 */
            {8'h00}, /* 0x6776 */
            {8'h00}, /* 0x6775 */
            {8'h00}, /* 0x6774 */
            {8'h00}, /* 0x6773 */
            {8'h00}, /* 0x6772 */
            {8'h00}, /* 0x6771 */
            {8'h00}, /* 0x6770 */
            {8'h00}, /* 0x676f */
            {8'h00}, /* 0x676e */
            {8'h00}, /* 0x676d */
            {8'h00}, /* 0x676c */
            {8'h00}, /* 0x676b */
            {8'h00}, /* 0x676a */
            {8'h00}, /* 0x6769 */
            {8'h00}, /* 0x6768 */
            {8'h00}, /* 0x6767 */
            {8'h00}, /* 0x6766 */
            {8'h00}, /* 0x6765 */
            {8'h00}, /* 0x6764 */
            {8'h00}, /* 0x6763 */
            {8'h00}, /* 0x6762 */
            {8'h00}, /* 0x6761 */
            {8'h00}, /* 0x6760 */
            {8'h00}, /* 0x675f */
            {8'h00}, /* 0x675e */
            {8'h00}, /* 0x675d */
            {8'h00}, /* 0x675c */
            {8'h00}, /* 0x675b */
            {8'h00}, /* 0x675a */
            {8'h00}, /* 0x6759 */
            {8'h00}, /* 0x6758 */
            {8'h00}, /* 0x6757 */
            {8'h00}, /* 0x6756 */
            {8'h00}, /* 0x6755 */
            {8'h00}, /* 0x6754 */
            {8'h00}, /* 0x6753 */
            {8'h00}, /* 0x6752 */
            {8'h00}, /* 0x6751 */
            {8'h00}, /* 0x6750 */
            {8'h00}, /* 0x674f */
            {8'h00}, /* 0x674e */
            {8'h00}, /* 0x674d */
            {8'h00}, /* 0x674c */
            {8'h00}, /* 0x674b */
            {8'h00}, /* 0x674a */
            {8'h00}, /* 0x6749 */
            {8'h00}, /* 0x6748 */
            {8'h00}, /* 0x6747 */
            {8'h00}, /* 0x6746 */
            {8'h00}, /* 0x6745 */
            {8'h00}, /* 0x6744 */
            {8'h00}, /* 0x6743 */
            {8'h00}, /* 0x6742 */
            {8'h00}, /* 0x6741 */
            {8'h00}, /* 0x6740 */
            {8'h00}, /* 0x673f */
            {8'h00}, /* 0x673e */
            {8'h00}, /* 0x673d */
            {8'h00}, /* 0x673c */
            {8'h00}, /* 0x673b */
            {8'h00}, /* 0x673a */
            {8'h00}, /* 0x6739 */
            {8'h00}, /* 0x6738 */
            {8'h00}, /* 0x6737 */
            {8'h00}, /* 0x6736 */
            {8'h00}, /* 0x6735 */
            {8'h00}, /* 0x6734 */
            {8'h00}, /* 0x6733 */
            {8'h00}, /* 0x6732 */
            {8'h00}, /* 0x6731 */
            {8'h00}, /* 0x6730 */
            {8'h00}, /* 0x672f */
            {8'h00}, /* 0x672e */
            {8'h00}, /* 0x672d */
            {8'h00}, /* 0x672c */
            {8'h00}, /* 0x672b */
            {8'h00}, /* 0x672a */
            {8'h00}, /* 0x6729 */
            {8'h00}, /* 0x6728 */
            {8'h00}, /* 0x6727 */
            {8'h00}, /* 0x6726 */
            {8'h00}, /* 0x6725 */
            {8'h00}, /* 0x6724 */
            {8'h00}, /* 0x6723 */
            {8'h00}, /* 0x6722 */
            {8'h00}, /* 0x6721 */
            {8'h00}, /* 0x6720 */
            {8'h00}, /* 0x671f */
            {8'h00}, /* 0x671e */
            {8'h00}, /* 0x671d */
            {8'h00}, /* 0x671c */
            {8'h00}, /* 0x671b */
            {8'h00}, /* 0x671a */
            {8'h00}, /* 0x6719 */
            {8'h00}, /* 0x6718 */
            {8'h00}, /* 0x6717 */
            {8'h00}, /* 0x6716 */
            {8'h00}, /* 0x6715 */
            {8'h00}, /* 0x6714 */
            {8'h00}, /* 0x6713 */
            {8'h00}, /* 0x6712 */
            {8'h00}, /* 0x6711 */
            {8'h00}, /* 0x6710 */
            {8'h00}, /* 0x670f */
            {8'h00}, /* 0x670e */
            {8'h00}, /* 0x670d */
            {8'h00}, /* 0x670c */
            {8'h00}, /* 0x670b */
            {8'h00}, /* 0x670a */
            {8'h00}, /* 0x6709 */
            {8'h00}, /* 0x6708 */
            {8'h00}, /* 0x6707 */
            {8'h00}, /* 0x6706 */
            {8'h00}, /* 0x6705 */
            {8'h00}, /* 0x6704 */
            {8'h00}, /* 0x6703 */
            {8'h00}, /* 0x6702 */
            {8'h00}, /* 0x6701 */
            {8'h00}, /* 0x6700 */
            {8'h00}, /* 0x66ff */
            {8'h00}, /* 0x66fe */
            {8'h00}, /* 0x66fd */
            {8'h00}, /* 0x66fc */
            {8'h00}, /* 0x66fb */
            {8'h00}, /* 0x66fa */
            {8'h00}, /* 0x66f9 */
            {8'h00}, /* 0x66f8 */
            {8'h00}, /* 0x66f7 */
            {8'h00}, /* 0x66f6 */
            {8'h00}, /* 0x66f5 */
            {8'h00}, /* 0x66f4 */
            {8'h00}, /* 0x66f3 */
            {8'h00}, /* 0x66f2 */
            {8'h00}, /* 0x66f1 */
            {8'h00}, /* 0x66f0 */
            {8'h00}, /* 0x66ef */
            {8'h00}, /* 0x66ee */
            {8'h00}, /* 0x66ed */
            {8'h00}, /* 0x66ec */
            {8'h00}, /* 0x66eb */
            {8'h00}, /* 0x66ea */
            {8'h00}, /* 0x66e9 */
            {8'h00}, /* 0x66e8 */
            {8'h00}, /* 0x66e7 */
            {8'h00}, /* 0x66e6 */
            {8'h00}, /* 0x66e5 */
            {8'h00}, /* 0x66e4 */
            {8'h00}, /* 0x66e3 */
            {8'h00}, /* 0x66e2 */
            {8'h00}, /* 0x66e1 */
            {8'h00}, /* 0x66e0 */
            {8'h00}, /* 0x66df */
            {8'h00}, /* 0x66de */
            {8'h00}, /* 0x66dd */
            {8'h00}, /* 0x66dc */
            {8'h00}, /* 0x66db */
            {8'h00}, /* 0x66da */
            {8'h00}, /* 0x66d9 */
            {8'h00}, /* 0x66d8 */
            {8'h00}, /* 0x66d7 */
            {8'h00}, /* 0x66d6 */
            {8'h00}, /* 0x66d5 */
            {8'h00}, /* 0x66d4 */
            {8'h00}, /* 0x66d3 */
            {8'h00}, /* 0x66d2 */
            {8'h00}, /* 0x66d1 */
            {8'h00}, /* 0x66d0 */
            {8'h00}, /* 0x66cf */
            {8'h00}, /* 0x66ce */
            {8'h00}, /* 0x66cd */
            {8'h00}, /* 0x66cc */
            {8'h00}, /* 0x66cb */
            {8'h00}, /* 0x66ca */
            {8'h00}, /* 0x66c9 */
            {8'h00}, /* 0x66c8 */
            {8'h00}, /* 0x66c7 */
            {8'h00}, /* 0x66c6 */
            {8'h00}, /* 0x66c5 */
            {8'h00}, /* 0x66c4 */
            {8'h00}, /* 0x66c3 */
            {8'h00}, /* 0x66c2 */
            {8'h00}, /* 0x66c1 */
            {8'h00}, /* 0x66c0 */
            {8'h00}, /* 0x66bf */
            {8'h00}, /* 0x66be */
            {8'h00}, /* 0x66bd */
            {8'h00}, /* 0x66bc */
            {8'h00}, /* 0x66bb */
            {8'h00}, /* 0x66ba */
            {8'h00}, /* 0x66b9 */
            {8'h00}, /* 0x66b8 */
            {8'h00}, /* 0x66b7 */
            {8'h00}, /* 0x66b6 */
            {8'h00}, /* 0x66b5 */
            {8'h00}, /* 0x66b4 */
            {8'h00}, /* 0x66b3 */
            {8'h00}, /* 0x66b2 */
            {8'h00}, /* 0x66b1 */
            {8'h00}, /* 0x66b0 */
            {8'h00}, /* 0x66af */
            {8'h00}, /* 0x66ae */
            {8'h00}, /* 0x66ad */
            {8'h00}, /* 0x66ac */
            {8'h00}, /* 0x66ab */
            {8'h00}, /* 0x66aa */
            {8'h00}, /* 0x66a9 */
            {8'h00}, /* 0x66a8 */
            {8'h00}, /* 0x66a7 */
            {8'h00}, /* 0x66a6 */
            {8'h00}, /* 0x66a5 */
            {8'h00}, /* 0x66a4 */
            {8'h00}, /* 0x66a3 */
            {8'h00}, /* 0x66a2 */
            {8'h00}, /* 0x66a1 */
            {8'h00}, /* 0x66a0 */
            {8'h00}, /* 0x669f */
            {8'h00}, /* 0x669e */
            {8'h00}, /* 0x669d */
            {8'h00}, /* 0x669c */
            {8'h00}, /* 0x669b */
            {8'h00}, /* 0x669a */
            {8'h00}, /* 0x6699 */
            {8'h00}, /* 0x6698 */
            {8'h00}, /* 0x6697 */
            {8'h00}, /* 0x6696 */
            {8'h00}, /* 0x6695 */
            {8'h00}, /* 0x6694 */
            {8'h00}, /* 0x6693 */
            {8'h00}, /* 0x6692 */
            {8'h00}, /* 0x6691 */
            {8'h00}, /* 0x6690 */
            {8'h00}, /* 0x668f */
            {8'h00}, /* 0x668e */
            {8'h00}, /* 0x668d */
            {8'h00}, /* 0x668c */
            {8'h00}, /* 0x668b */
            {8'h00}, /* 0x668a */
            {8'h00}, /* 0x6689 */
            {8'h00}, /* 0x6688 */
            {8'h00}, /* 0x6687 */
            {8'h00}, /* 0x6686 */
            {8'h00}, /* 0x6685 */
            {8'h00}, /* 0x6684 */
            {8'h00}, /* 0x6683 */
            {8'h00}, /* 0x6682 */
            {8'h00}, /* 0x6681 */
            {8'h00}, /* 0x6680 */
            {8'h00}, /* 0x667f */
            {8'h00}, /* 0x667e */
            {8'h00}, /* 0x667d */
            {8'h00}, /* 0x667c */
            {8'h00}, /* 0x667b */
            {8'h00}, /* 0x667a */
            {8'h00}, /* 0x6679 */
            {8'h00}, /* 0x6678 */
            {8'h00}, /* 0x6677 */
            {8'h00}, /* 0x6676 */
            {8'h00}, /* 0x6675 */
            {8'h00}, /* 0x6674 */
            {8'h00}, /* 0x6673 */
            {8'h00}, /* 0x6672 */
            {8'h00}, /* 0x6671 */
            {8'h00}, /* 0x6670 */
            {8'h00}, /* 0x666f */
            {8'h00}, /* 0x666e */
            {8'h00}, /* 0x666d */
            {8'h00}, /* 0x666c */
            {8'h00}, /* 0x666b */
            {8'h00}, /* 0x666a */
            {8'h00}, /* 0x6669 */
            {8'h00}, /* 0x6668 */
            {8'h00}, /* 0x6667 */
            {8'h00}, /* 0x6666 */
            {8'h00}, /* 0x6665 */
            {8'h00}, /* 0x6664 */
            {8'h00}, /* 0x6663 */
            {8'h00}, /* 0x6662 */
            {8'h00}, /* 0x6661 */
            {8'h00}, /* 0x6660 */
            {8'h00}, /* 0x665f */
            {8'h00}, /* 0x665e */
            {8'h00}, /* 0x665d */
            {8'h00}, /* 0x665c */
            {8'h00}, /* 0x665b */
            {8'h00}, /* 0x665a */
            {8'h00}, /* 0x6659 */
            {8'h00}, /* 0x6658 */
            {8'h00}, /* 0x6657 */
            {8'h00}, /* 0x6656 */
            {8'h00}, /* 0x6655 */
            {8'h00}, /* 0x6654 */
            {8'h00}, /* 0x6653 */
            {8'h00}, /* 0x6652 */
            {8'h00}, /* 0x6651 */
            {8'h00}, /* 0x6650 */
            {8'h00}, /* 0x664f */
            {8'h00}, /* 0x664e */
            {8'h00}, /* 0x664d */
            {8'h00}, /* 0x664c */
            {8'h00}, /* 0x664b */
            {8'h00}, /* 0x664a */
            {8'h00}, /* 0x6649 */
            {8'h00}, /* 0x6648 */
            {8'h00}, /* 0x6647 */
            {8'h00}, /* 0x6646 */
            {8'h00}, /* 0x6645 */
            {8'h00}, /* 0x6644 */
            {8'h00}, /* 0x6643 */
            {8'h00}, /* 0x6642 */
            {8'h00}, /* 0x6641 */
            {8'h00}, /* 0x6640 */
            {8'h00}, /* 0x663f */
            {8'h00}, /* 0x663e */
            {8'h00}, /* 0x663d */
            {8'h00}, /* 0x663c */
            {8'h00}, /* 0x663b */
            {8'h00}, /* 0x663a */
            {8'h00}, /* 0x6639 */
            {8'h00}, /* 0x6638 */
            {8'h00}, /* 0x6637 */
            {8'h00}, /* 0x6636 */
            {8'h00}, /* 0x6635 */
            {8'h00}, /* 0x6634 */
            {8'h00}, /* 0x6633 */
            {8'h00}, /* 0x6632 */
            {8'h00}, /* 0x6631 */
            {8'h00}, /* 0x6630 */
            {8'h00}, /* 0x662f */
            {8'h00}, /* 0x662e */
            {8'h00}, /* 0x662d */
            {8'h00}, /* 0x662c */
            {8'h00}, /* 0x662b */
            {8'h00}, /* 0x662a */
            {8'h00}, /* 0x6629 */
            {8'h00}, /* 0x6628 */
            {8'h00}, /* 0x6627 */
            {8'h00}, /* 0x6626 */
            {8'h00}, /* 0x6625 */
            {8'h00}, /* 0x6624 */
            {8'h00}, /* 0x6623 */
            {8'h00}, /* 0x6622 */
            {8'h00}, /* 0x6621 */
            {8'h00}, /* 0x6620 */
            {8'h00}, /* 0x661f */
            {8'h00}, /* 0x661e */
            {8'h00}, /* 0x661d */
            {8'h00}, /* 0x661c */
            {8'h00}, /* 0x661b */
            {8'h00}, /* 0x661a */
            {8'h00}, /* 0x6619 */
            {8'h00}, /* 0x6618 */
            {8'h00}, /* 0x6617 */
            {8'h00}, /* 0x6616 */
            {8'h00}, /* 0x6615 */
            {8'h00}, /* 0x6614 */
            {8'h00}, /* 0x6613 */
            {8'h00}, /* 0x6612 */
            {8'h00}, /* 0x6611 */
            {8'h00}, /* 0x6610 */
            {8'h00}, /* 0x660f */
            {8'h00}, /* 0x660e */
            {8'h00}, /* 0x660d */
            {8'h00}, /* 0x660c */
            {8'h00}, /* 0x660b */
            {8'h00}, /* 0x660a */
            {8'h00}, /* 0x6609 */
            {8'h00}, /* 0x6608 */
            {8'h00}, /* 0x6607 */
            {8'h00}, /* 0x6606 */
            {8'h00}, /* 0x6605 */
            {8'h00}, /* 0x6604 */
            {8'h00}, /* 0x6603 */
            {8'h00}, /* 0x6602 */
            {8'h00}, /* 0x6601 */
            {8'h00}, /* 0x6600 */
            {8'h00}, /* 0x65ff */
            {8'h00}, /* 0x65fe */
            {8'h00}, /* 0x65fd */
            {8'h00}, /* 0x65fc */
            {8'h00}, /* 0x65fb */
            {8'h00}, /* 0x65fa */
            {8'h00}, /* 0x65f9 */
            {8'h00}, /* 0x65f8 */
            {8'h00}, /* 0x65f7 */
            {8'h00}, /* 0x65f6 */
            {8'h00}, /* 0x65f5 */
            {8'h00}, /* 0x65f4 */
            {8'h00}, /* 0x65f3 */
            {8'h00}, /* 0x65f2 */
            {8'h00}, /* 0x65f1 */
            {8'h00}, /* 0x65f0 */
            {8'h00}, /* 0x65ef */
            {8'h00}, /* 0x65ee */
            {8'h00}, /* 0x65ed */
            {8'h00}, /* 0x65ec */
            {8'h00}, /* 0x65eb */
            {8'h00}, /* 0x65ea */
            {8'h00}, /* 0x65e9 */
            {8'h00}, /* 0x65e8 */
            {8'h00}, /* 0x65e7 */
            {8'h00}, /* 0x65e6 */
            {8'h00}, /* 0x65e5 */
            {8'h00}, /* 0x65e4 */
            {8'h00}, /* 0x65e3 */
            {8'h00}, /* 0x65e2 */
            {8'h00}, /* 0x65e1 */
            {8'h00}, /* 0x65e0 */
            {8'h00}, /* 0x65df */
            {8'h00}, /* 0x65de */
            {8'h00}, /* 0x65dd */
            {8'h00}, /* 0x65dc */
            {8'h00}, /* 0x65db */
            {8'h00}, /* 0x65da */
            {8'h00}, /* 0x65d9 */
            {8'h00}, /* 0x65d8 */
            {8'h00}, /* 0x65d7 */
            {8'h00}, /* 0x65d6 */
            {8'h00}, /* 0x65d5 */
            {8'h00}, /* 0x65d4 */
            {8'h00}, /* 0x65d3 */
            {8'h00}, /* 0x65d2 */
            {8'h00}, /* 0x65d1 */
            {8'h00}, /* 0x65d0 */
            {8'h00}, /* 0x65cf */
            {8'h00}, /* 0x65ce */
            {8'h00}, /* 0x65cd */
            {8'h00}, /* 0x65cc */
            {8'h00}, /* 0x65cb */
            {8'h00}, /* 0x65ca */
            {8'h00}, /* 0x65c9 */
            {8'h00}, /* 0x65c8 */
            {8'h00}, /* 0x65c7 */
            {8'h00}, /* 0x65c6 */
            {8'h00}, /* 0x65c5 */
            {8'h00}, /* 0x65c4 */
            {8'h00}, /* 0x65c3 */
            {8'h00}, /* 0x65c2 */
            {8'h00}, /* 0x65c1 */
            {8'h00}, /* 0x65c0 */
            {8'h00}, /* 0x65bf */
            {8'h00}, /* 0x65be */
            {8'h00}, /* 0x65bd */
            {8'h00}, /* 0x65bc */
            {8'h00}, /* 0x65bb */
            {8'h00}, /* 0x65ba */
            {8'h00}, /* 0x65b9 */
            {8'h00}, /* 0x65b8 */
            {8'h00}, /* 0x65b7 */
            {8'h00}, /* 0x65b6 */
            {8'h00}, /* 0x65b5 */
            {8'h00}, /* 0x65b4 */
            {8'h00}, /* 0x65b3 */
            {8'h00}, /* 0x65b2 */
            {8'h00}, /* 0x65b1 */
            {8'h00}, /* 0x65b0 */
            {8'h00}, /* 0x65af */
            {8'h00}, /* 0x65ae */
            {8'h00}, /* 0x65ad */
            {8'h00}, /* 0x65ac */
            {8'h00}, /* 0x65ab */
            {8'h00}, /* 0x65aa */
            {8'h00}, /* 0x65a9 */
            {8'h00}, /* 0x65a8 */
            {8'h00}, /* 0x65a7 */
            {8'h00}, /* 0x65a6 */
            {8'h00}, /* 0x65a5 */
            {8'h00}, /* 0x65a4 */
            {8'h00}, /* 0x65a3 */
            {8'h00}, /* 0x65a2 */
            {8'h00}, /* 0x65a1 */
            {8'h00}, /* 0x65a0 */
            {8'h00}, /* 0x659f */
            {8'h00}, /* 0x659e */
            {8'h00}, /* 0x659d */
            {8'h00}, /* 0x659c */
            {8'h00}, /* 0x659b */
            {8'h00}, /* 0x659a */
            {8'h00}, /* 0x6599 */
            {8'h00}, /* 0x6598 */
            {8'h00}, /* 0x6597 */
            {8'h00}, /* 0x6596 */
            {8'h00}, /* 0x6595 */
            {8'h00}, /* 0x6594 */
            {8'h00}, /* 0x6593 */
            {8'h00}, /* 0x6592 */
            {8'h00}, /* 0x6591 */
            {8'h00}, /* 0x6590 */
            {8'h00}, /* 0x658f */
            {8'h00}, /* 0x658e */
            {8'h00}, /* 0x658d */
            {8'h00}, /* 0x658c */
            {8'h00}, /* 0x658b */
            {8'h00}, /* 0x658a */
            {8'h00}, /* 0x6589 */
            {8'h00}, /* 0x6588 */
            {8'h00}, /* 0x6587 */
            {8'h00}, /* 0x6586 */
            {8'h00}, /* 0x6585 */
            {8'h00}, /* 0x6584 */
            {8'h00}, /* 0x6583 */
            {8'h00}, /* 0x6582 */
            {8'h00}, /* 0x6581 */
            {8'h00}, /* 0x6580 */
            {8'h00}, /* 0x657f */
            {8'h00}, /* 0x657e */
            {8'h00}, /* 0x657d */
            {8'h00}, /* 0x657c */
            {8'h00}, /* 0x657b */
            {8'h00}, /* 0x657a */
            {8'h00}, /* 0x6579 */
            {8'h00}, /* 0x6578 */
            {8'h00}, /* 0x6577 */
            {8'h00}, /* 0x6576 */
            {8'h00}, /* 0x6575 */
            {8'h00}, /* 0x6574 */
            {8'h00}, /* 0x6573 */
            {8'h00}, /* 0x6572 */
            {8'h00}, /* 0x6571 */
            {8'h00}, /* 0x6570 */
            {8'h00}, /* 0x656f */
            {8'h00}, /* 0x656e */
            {8'h00}, /* 0x656d */
            {8'h00}, /* 0x656c */
            {8'h00}, /* 0x656b */
            {8'h00}, /* 0x656a */
            {8'h00}, /* 0x6569 */
            {8'h00}, /* 0x6568 */
            {8'h00}, /* 0x6567 */
            {8'h00}, /* 0x6566 */
            {8'h00}, /* 0x6565 */
            {8'h00}, /* 0x6564 */
            {8'h00}, /* 0x6563 */
            {8'h00}, /* 0x6562 */
            {8'h00}, /* 0x6561 */
            {8'h00}, /* 0x6560 */
            {8'h00}, /* 0x655f */
            {8'h00}, /* 0x655e */
            {8'h00}, /* 0x655d */
            {8'h00}, /* 0x655c */
            {8'h00}, /* 0x655b */
            {8'h00}, /* 0x655a */
            {8'h00}, /* 0x6559 */
            {8'h00}, /* 0x6558 */
            {8'h00}, /* 0x6557 */
            {8'h00}, /* 0x6556 */
            {8'h00}, /* 0x6555 */
            {8'h00}, /* 0x6554 */
            {8'h00}, /* 0x6553 */
            {8'h00}, /* 0x6552 */
            {8'h00}, /* 0x6551 */
            {8'h00}, /* 0x6550 */
            {8'h00}, /* 0x654f */
            {8'h00}, /* 0x654e */
            {8'h00}, /* 0x654d */
            {8'h00}, /* 0x654c */
            {8'h00}, /* 0x654b */
            {8'h00}, /* 0x654a */
            {8'h00}, /* 0x6549 */
            {8'h00}, /* 0x6548 */
            {8'h00}, /* 0x6547 */
            {8'h00}, /* 0x6546 */
            {8'h00}, /* 0x6545 */
            {8'h00}, /* 0x6544 */
            {8'h00}, /* 0x6543 */
            {8'h00}, /* 0x6542 */
            {8'h00}, /* 0x6541 */
            {8'h00}, /* 0x6540 */
            {8'h00}, /* 0x653f */
            {8'h00}, /* 0x653e */
            {8'h00}, /* 0x653d */
            {8'h00}, /* 0x653c */
            {8'h00}, /* 0x653b */
            {8'h00}, /* 0x653a */
            {8'h00}, /* 0x6539 */
            {8'h00}, /* 0x6538 */
            {8'h00}, /* 0x6537 */
            {8'h00}, /* 0x6536 */
            {8'h00}, /* 0x6535 */
            {8'h00}, /* 0x6534 */
            {8'h00}, /* 0x6533 */
            {8'h00}, /* 0x6532 */
            {8'h00}, /* 0x6531 */
            {8'h00}, /* 0x6530 */
            {8'h00}, /* 0x652f */
            {8'h00}, /* 0x652e */
            {8'h00}, /* 0x652d */
            {8'h00}, /* 0x652c */
            {8'h00}, /* 0x652b */
            {8'h00}, /* 0x652a */
            {8'h00}, /* 0x6529 */
            {8'h00}, /* 0x6528 */
            {8'h00}, /* 0x6527 */
            {8'h00}, /* 0x6526 */
            {8'h00}, /* 0x6525 */
            {8'h00}, /* 0x6524 */
            {8'h00}, /* 0x6523 */
            {8'h00}, /* 0x6522 */
            {8'h00}, /* 0x6521 */
            {8'h00}, /* 0x6520 */
            {8'h00}, /* 0x651f */
            {8'h00}, /* 0x651e */
            {8'h00}, /* 0x651d */
            {8'h00}, /* 0x651c */
            {8'h00}, /* 0x651b */
            {8'h00}, /* 0x651a */
            {8'h00}, /* 0x6519 */
            {8'h00}, /* 0x6518 */
            {8'h00}, /* 0x6517 */
            {8'h00}, /* 0x6516 */
            {8'h00}, /* 0x6515 */
            {8'h00}, /* 0x6514 */
            {8'h00}, /* 0x6513 */
            {8'h00}, /* 0x6512 */
            {8'h00}, /* 0x6511 */
            {8'h00}, /* 0x6510 */
            {8'h00}, /* 0x650f */
            {8'h00}, /* 0x650e */
            {8'h00}, /* 0x650d */
            {8'h00}, /* 0x650c */
            {8'h00}, /* 0x650b */
            {8'h00}, /* 0x650a */
            {8'h00}, /* 0x6509 */
            {8'h00}, /* 0x6508 */
            {8'h00}, /* 0x6507 */
            {8'h00}, /* 0x6506 */
            {8'h00}, /* 0x6505 */
            {8'h00}, /* 0x6504 */
            {8'h00}, /* 0x6503 */
            {8'h00}, /* 0x6502 */
            {8'h00}, /* 0x6501 */
            {8'h00}, /* 0x6500 */
            {8'h00}, /* 0x64ff */
            {8'h00}, /* 0x64fe */
            {8'h00}, /* 0x64fd */
            {8'h00}, /* 0x64fc */
            {8'h00}, /* 0x64fb */
            {8'h00}, /* 0x64fa */
            {8'h00}, /* 0x64f9 */
            {8'h00}, /* 0x64f8 */
            {8'h00}, /* 0x64f7 */
            {8'h00}, /* 0x64f6 */
            {8'h00}, /* 0x64f5 */
            {8'h00}, /* 0x64f4 */
            {8'h00}, /* 0x64f3 */
            {8'h00}, /* 0x64f2 */
            {8'h00}, /* 0x64f1 */
            {8'h00}, /* 0x64f0 */
            {8'h00}, /* 0x64ef */
            {8'h00}, /* 0x64ee */
            {8'h00}, /* 0x64ed */
            {8'h00}, /* 0x64ec */
            {8'h00}, /* 0x64eb */
            {8'h00}, /* 0x64ea */
            {8'h00}, /* 0x64e9 */
            {8'h00}, /* 0x64e8 */
            {8'h00}, /* 0x64e7 */
            {8'h00}, /* 0x64e6 */
            {8'h00}, /* 0x64e5 */
            {8'h00}, /* 0x64e4 */
            {8'h00}, /* 0x64e3 */
            {8'h00}, /* 0x64e2 */
            {8'h00}, /* 0x64e1 */
            {8'h00}, /* 0x64e0 */
            {8'h00}, /* 0x64df */
            {8'h00}, /* 0x64de */
            {8'h00}, /* 0x64dd */
            {8'h00}, /* 0x64dc */
            {8'h00}, /* 0x64db */
            {8'h00}, /* 0x64da */
            {8'h00}, /* 0x64d9 */
            {8'h00}, /* 0x64d8 */
            {8'h00}, /* 0x64d7 */
            {8'h00}, /* 0x64d6 */
            {8'h00}, /* 0x64d5 */
            {8'h00}, /* 0x64d4 */
            {8'h00}, /* 0x64d3 */
            {8'h00}, /* 0x64d2 */
            {8'h00}, /* 0x64d1 */
            {8'h00}, /* 0x64d0 */
            {8'h00}, /* 0x64cf */
            {8'h00}, /* 0x64ce */
            {8'h00}, /* 0x64cd */
            {8'h00}, /* 0x64cc */
            {8'h00}, /* 0x64cb */
            {8'h00}, /* 0x64ca */
            {8'h00}, /* 0x64c9 */
            {8'h00}, /* 0x64c8 */
            {8'h00}, /* 0x64c7 */
            {8'h00}, /* 0x64c6 */
            {8'h00}, /* 0x64c5 */
            {8'h00}, /* 0x64c4 */
            {8'h00}, /* 0x64c3 */
            {8'h00}, /* 0x64c2 */
            {8'h00}, /* 0x64c1 */
            {8'h00}, /* 0x64c0 */
            {8'h00}, /* 0x64bf */
            {8'h00}, /* 0x64be */
            {8'h00}, /* 0x64bd */
            {8'h00}, /* 0x64bc */
            {8'h00}, /* 0x64bb */
            {8'h00}, /* 0x64ba */
            {8'h00}, /* 0x64b9 */
            {8'h00}, /* 0x64b8 */
            {8'h00}, /* 0x64b7 */
            {8'h00}, /* 0x64b6 */
            {8'h00}, /* 0x64b5 */
            {8'h00}, /* 0x64b4 */
            {8'h00}, /* 0x64b3 */
            {8'h00}, /* 0x64b2 */
            {8'h00}, /* 0x64b1 */
            {8'h00}, /* 0x64b0 */
            {8'h00}, /* 0x64af */
            {8'h00}, /* 0x64ae */
            {8'h00}, /* 0x64ad */
            {8'h00}, /* 0x64ac */
            {8'h00}, /* 0x64ab */
            {8'h00}, /* 0x64aa */
            {8'h00}, /* 0x64a9 */
            {8'h00}, /* 0x64a8 */
            {8'h00}, /* 0x64a7 */
            {8'h00}, /* 0x64a6 */
            {8'h00}, /* 0x64a5 */
            {8'h00}, /* 0x64a4 */
            {8'h00}, /* 0x64a3 */
            {8'h00}, /* 0x64a2 */
            {8'h00}, /* 0x64a1 */
            {8'h00}, /* 0x64a0 */
            {8'h00}, /* 0x649f */
            {8'h00}, /* 0x649e */
            {8'h00}, /* 0x649d */
            {8'h00}, /* 0x649c */
            {8'h00}, /* 0x649b */
            {8'h00}, /* 0x649a */
            {8'h00}, /* 0x6499 */
            {8'h00}, /* 0x6498 */
            {8'h00}, /* 0x6497 */
            {8'h00}, /* 0x6496 */
            {8'h00}, /* 0x6495 */
            {8'h00}, /* 0x6494 */
            {8'h00}, /* 0x6493 */
            {8'h00}, /* 0x6492 */
            {8'h00}, /* 0x6491 */
            {8'h00}, /* 0x6490 */
            {8'h00}, /* 0x648f */
            {8'h00}, /* 0x648e */
            {8'h00}, /* 0x648d */
            {8'h00}, /* 0x648c */
            {8'h00}, /* 0x648b */
            {8'h00}, /* 0x648a */
            {8'h00}, /* 0x6489 */
            {8'h00}, /* 0x6488 */
            {8'h00}, /* 0x6487 */
            {8'h00}, /* 0x6486 */
            {8'h00}, /* 0x6485 */
            {8'h00}, /* 0x6484 */
            {8'h00}, /* 0x6483 */
            {8'h00}, /* 0x6482 */
            {8'h00}, /* 0x6481 */
            {8'h00}, /* 0x6480 */
            {8'h00}, /* 0x647f */
            {8'h00}, /* 0x647e */
            {8'h00}, /* 0x647d */
            {8'h00}, /* 0x647c */
            {8'h00}, /* 0x647b */
            {8'h00}, /* 0x647a */
            {8'h00}, /* 0x6479 */
            {8'h00}, /* 0x6478 */
            {8'h00}, /* 0x6477 */
            {8'h00}, /* 0x6476 */
            {8'h00}, /* 0x6475 */
            {8'h00}, /* 0x6474 */
            {8'h00}, /* 0x6473 */
            {8'h00}, /* 0x6472 */
            {8'h00}, /* 0x6471 */
            {8'h00}, /* 0x6470 */
            {8'h00}, /* 0x646f */
            {8'h00}, /* 0x646e */
            {8'h00}, /* 0x646d */
            {8'h00}, /* 0x646c */
            {8'h00}, /* 0x646b */
            {8'h00}, /* 0x646a */
            {8'h00}, /* 0x6469 */
            {8'h00}, /* 0x6468 */
            {8'h00}, /* 0x6467 */
            {8'h00}, /* 0x6466 */
            {8'h00}, /* 0x6465 */
            {8'h00}, /* 0x6464 */
            {8'h00}, /* 0x6463 */
            {8'h00}, /* 0x6462 */
            {8'h00}, /* 0x6461 */
            {8'h00}, /* 0x6460 */
            {8'h00}, /* 0x645f */
            {8'h00}, /* 0x645e */
            {8'h00}, /* 0x645d */
            {8'h00}, /* 0x645c */
            {8'h00}, /* 0x645b */
            {8'h00}, /* 0x645a */
            {8'h00}, /* 0x6459 */
            {8'h00}, /* 0x6458 */
            {8'h00}, /* 0x6457 */
            {8'h00}, /* 0x6456 */
            {8'h00}, /* 0x6455 */
            {8'h00}, /* 0x6454 */
            {8'h00}, /* 0x6453 */
            {8'h00}, /* 0x6452 */
            {8'h00}, /* 0x6451 */
            {8'h00}, /* 0x6450 */
            {8'h00}, /* 0x644f */
            {8'h00}, /* 0x644e */
            {8'h00}, /* 0x644d */
            {8'h00}, /* 0x644c */
            {8'h00}, /* 0x644b */
            {8'h00}, /* 0x644a */
            {8'h00}, /* 0x6449 */
            {8'h00}, /* 0x6448 */
            {8'h00}, /* 0x6447 */
            {8'h00}, /* 0x6446 */
            {8'h00}, /* 0x6445 */
            {8'h00}, /* 0x6444 */
            {8'h00}, /* 0x6443 */
            {8'h00}, /* 0x6442 */
            {8'h00}, /* 0x6441 */
            {8'h00}, /* 0x6440 */
            {8'h00}, /* 0x643f */
            {8'h00}, /* 0x643e */
            {8'h00}, /* 0x643d */
            {8'h00}, /* 0x643c */
            {8'h00}, /* 0x643b */
            {8'h00}, /* 0x643a */
            {8'h00}, /* 0x6439 */
            {8'h00}, /* 0x6438 */
            {8'h00}, /* 0x6437 */
            {8'h00}, /* 0x6436 */
            {8'h00}, /* 0x6435 */
            {8'h00}, /* 0x6434 */
            {8'h00}, /* 0x6433 */
            {8'h00}, /* 0x6432 */
            {8'h00}, /* 0x6431 */
            {8'h00}, /* 0x6430 */
            {8'h00}, /* 0x642f */
            {8'h00}, /* 0x642e */
            {8'h00}, /* 0x642d */
            {8'h00}, /* 0x642c */
            {8'h00}, /* 0x642b */
            {8'h00}, /* 0x642a */
            {8'h00}, /* 0x6429 */
            {8'h00}, /* 0x6428 */
            {8'h00}, /* 0x6427 */
            {8'h00}, /* 0x6426 */
            {8'h00}, /* 0x6425 */
            {8'h00}, /* 0x6424 */
            {8'h00}, /* 0x6423 */
            {8'h00}, /* 0x6422 */
            {8'h00}, /* 0x6421 */
            {8'h00}, /* 0x6420 */
            {8'h00}, /* 0x641f */
            {8'h00}, /* 0x641e */
            {8'h00}, /* 0x641d */
            {8'h00}, /* 0x641c */
            {8'h00}, /* 0x641b */
            {8'h00}, /* 0x641a */
            {8'h00}, /* 0x6419 */
            {8'h00}, /* 0x6418 */
            {8'h00}, /* 0x6417 */
            {8'h00}, /* 0x6416 */
            {8'h00}, /* 0x6415 */
            {8'h00}, /* 0x6414 */
            {8'h00}, /* 0x6413 */
            {8'h00}, /* 0x6412 */
            {8'h00}, /* 0x6411 */
            {8'h00}, /* 0x6410 */
            {8'h00}, /* 0x640f */
            {8'h00}, /* 0x640e */
            {8'h00}, /* 0x640d */
            {8'h00}, /* 0x640c */
            {8'h00}, /* 0x640b */
            {8'h00}, /* 0x640a */
            {8'h00}, /* 0x6409 */
            {8'h00}, /* 0x6408 */
            {8'h00}, /* 0x6407 */
            {8'h00}, /* 0x6406 */
            {8'h00}, /* 0x6405 */
            {8'h00}, /* 0x6404 */
            {8'h00}, /* 0x6403 */
            {8'h00}, /* 0x6402 */
            {8'h00}, /* 0x6401 */
            {8'h00}, /* 0x6400 */
            {8'h00}, /* 0x63ff */
            {8'h00}, /* 0x63fe */
            {8'h00}, /* 0x63fd */
            {8'h00}, /* 0x63fc */
            {8'h00}, /* 0x63fb */
            {8'h00}, /* 0x63fa */
            {8'h00}, /* 0x63f9 */
            {8'h00}, /* 0x63f8 */
            {8'h00}, /* 0x63f7 */
            {8'h00}, /* 0x63f6 */
            {8'h00}, /* 0x63f5 */
            {8'h00}, /* 0x63f4 */
            {8'h00}, /* 0x63f3 */
            {8'h00}, /* 0x63f2 */
            {8'h00}, /* 0x63f1 */
            {8'h00}, /* 0x63f0 */
            {8'h00}, /* 0x63ef */
            {8'h00}, /* 0x63ee */
            {8'h00}, /* 0x63ed */
            {8'h00}, /* 0x63ec */
            {8'h00}, /* 0x63eb */
            {8'h00}, /* 0x63ea */
            {8'h00}, /* 0x63e9 */
            {8'h00}, /* 0x63e8 */
            {8'h00}, /* 0x63e7 */
            {8'h00}, /* 0x63e6 */
            {8'h00}, /* 0x63e5 */
            {8'h00}, /* 0x63e4 */
            {8'h00}, /* 0x63e3 */
            {8'h00}, /* 0x63e2 */
            {8'h00}, /* 0x63e1 */
            {8'h00}, /* 0x63e0 */
            {8'h00}, /* 0x63df */
            {8'h00}, /* 0x63de */
            {8'h00}, /* 0x63dd */
            {8'h00}, /* 0x63dc */
            {8'h00}, /* 0x63db */
            {8'h00}, /* 0x63da */
            {8'h00}, /* 0x63d9 */
            {8'h00}, /* 0x63d8 */
            {8'h00}, /* 0x63d7 */
            {8'h00}, /* 0x63d6 */
            {8'h00}, /* 0x63d5 */
            {8'h00}, /* 0x63d4 */
            {8'h00}, /* 0x63d3 */
            {8'h00}, /* 0x63d2 */
            {8'h00}, /* 0x63d1 */
            {8'h00}, /* 0x63d0 */
            {8'h00}, /* 0x63cf */
            {8'h00}, /* 0x63ce */
            {8'h00}, /* 0x63cd */
            {8'h00}, /* 0x63cc */
            {8'h00}, /* 0x63cb */
            {8'h00}, /* 0x63ca */
            {8'h00}, /* 0x63c9 */
            {8'h00}, /* 0x63c8 */
            {8'h00}, /* 0x63c7 */
            {8'h00}, /* 0x63c6 */
            {8'h00}, /* 0x63c5 */
            {8'h00}, /* 0x63c4 */
            {8'h00}, /* 0x63c3 */
            {8'h00}, /* 0x63c2 */
            {8'h00}, /* 0x63c1 */
            {8'h00}, /* 0x63c0 */
            {8'h00}, /* 0x63bf */
            {8'h00}, /* 0x63be */
            {8'h00}, /* 0x63bd */
            {8'h00}, /* 0x63bc */
            {8'h00}, /* 0x63bb */
            {8'h00}, /* 0x63ba */
            {8'h00}, /* 0x63b9 */
            {8'h00}, /* 0x63b8 */
            {8'h00}, /* 0x63b7 */
            {8'h00}, /* 0x63b6 */
            {8'h00}, /* 0x63b5 */
            {8'h00}, /* 0x63b4 */
            {8'h00}, /* 0x63b3 */
            {8'h00}, /* 0x63b2 */
            {8'h00}, /* 0x63b1 */
            {8'h00}, /* 0x63b0 */
            {8'h00}, /* 0x63af */
            {8'h00}, /* 0x63ae */
            {8'h00}, /* 0x63ad */
            {8'h00}, /* 0x63ac */
            {8'h00}, /* 0x63ab */
            {8'h00}, /* 0x63aa */
            {8'h00}, /* 0x63a9 */
            {8'h00}, /* 0x63a8 */
            {8'h00}, /* 0x63a7 */
            {8'h00}, /* 0x63a6 */
            {8'h00}, /* 0x63a5 */
            {8'h00}, /* 0x63a4 */
            {8'h00}, /* 0x63a3 */
            {8'h00}, /* 0x63a2 */
            {8'h00}, /* 0x63a1 */
            {8'h00}, /* 0x63a0 */
            {8'h00}, /* 0x639f */
            {8'h00}, /* 0x639e */
            {8'h00}, /* 0x639d */
            {8'h00}, /* 0x639c */
            {8'h00}, /* 0x639b */
            {8'h00}, /* 0x639a */
            {8'h00}, /* 0x6399 */
            {8'h00}, /* 0x6398 */
            {8'h00}, /* 0x6397 */
            {8'h00}, /* 0x6396 */
            {8'h00}, /* 0x6395 */
            {8'h00}, /* 0x6394 */
            {8'h00}, /* 0x6393 */
            {8'h00}, /* 0x6392 */
            {8'h00}, /* 0x6391 */
            {8'h00}, /* 0x6390 */
            {8'h00}, /* 0x638f */
            {8'h00}, /* 0x638e */
            {8'h00}, /* 0x638d */
            {8'h00}, /* 0x638c */
            {8'h00}, /* 0x638b */
            {8'h00}, /* 0x638a */
            {8'h00}, /* 0x6389 */
            {8'h00}, /* 0x6388 */
            {8'h00}, /* 0x6387 */
            {8'h00}, /* 0x6386 */
            {8'h00}, /* 0x6385 */
            {8'h00}, /* 0x6384 */
            {8'h00}, /* 0x6383 */
            {8'h00}, /* 0x6382 */
            {8'h00}, /* 0x6381 */
            {8'h00}, /* 0x6380 */
            {8'h00}, /* 0x637f */
            {8'h00}, /* 0x637e */
            {8'h00}, /* 0x637d */
            {8'h00}, /* 0x637c */
            {8'h00}, /* 0x637b */
            {8'h00}, /* 0x637a */
            {8'h00}, /* 0x6379 */
            {8'h00}, /* 0x6378 */
            {8'h00}, /* 0x6377 */
            {8'h00}, /* 0x6376 */
            {8'h00}, /* 0x6375 */
            {8'h00}, /* 0x6374 */
            {8'h00}, /* 0x6373 */
            {8'h00}, /* 0x6372 */
            {8'h00}, /* 0x6371 */
            {8'h00}, /* 0x6370 */
            {8'h00}, /* 0x636f */
            {8'h00}, /* 0x636e */
            {8'h00}, /* 0x636d */
            {8'h00}, /* 0x636c */
            {8'h00}, /* 0x636b */
            {8'h00}, /* 0x636a */
            {8'h00}, /* 0x6369 */
            {8'h00}, /* 0x6368 */
            {8'h00}, /* 0x6367 */
            {8'h00}, /* 0x6366 */
            {8'h00}, /* 0x6365 */
            {8'h00}, /* 0x6364 */
            {8'h00}, /* 0x6363 */
            {8'h00}, /* 0x6362 */
            {8'h00}, /* 0x6361 */
            {8'h00}, /* 0x6360 */
            {8'h00}, /* 0x635f */
            {8'h00}, /* 0x635e */
            {8'h00}, /* 0x635d */
            {8'h00}, /* 0x635c */
            {8'h00}, /* 0x635b */
            {8'h00}, /* 0x635a */
            {8'h00}, /* 0x6359 */
            {8'h00}, /* 0x6358 */
            {8'h00}, /* 0x6357 */
            {8'h00}, /* 0x6356 */
            {8'h00}, /* 0x6355 */
            {8'h00}, /* 0x6354 */
            {8'h00}, /* 0x6353 */
            {8'h00}, /* 0x6352 */
            {8'h00}, /* 0x6351 */
            {8'h00}, /* 0x6350 */
            {8'h00}, /* 0x634f */
            {8'h00}, /* 0x634e */
            {8'h00}, /* 0x634d */
            {8'h00}, /* 0x634c */
            {8'h00}, /* 0x634b */
            {8'h00}, /* 0x634a */
            {8'h00}, /* 0x6349 */
            {8'h00}, /* 0x6348 */
            {8'h00}, /* 0x6347 */
            {8'h00}, /* 0x6346 */
            {8'h00}, /* 0x6345 */
            {8'h00}, /* 0x6344 */
            {8'h00}, /* 0x6343 */
            {8'h00}, /* 0x6342 */
            {8'h00}, /* 0x6341 */
            {8'h00}, /* 0x6340 */
            {8'h00}, /* 0x633f */
            {8'h00}, /* 0x633e */
            {8'h00}, /* 0x633d */
            {8'h00}, /* 0x633c */
            {8'h00}, /* 0x633b */
            {8'h00}, /* 0x633a */
            {8'h00}, /* 0x6339 */
            {8'h00}, /* 0x6338 */
            {8'h00}, /* 0x6337 */
            {8'h00}, /* 0x6336 */
            {8'h00}, /* 0x6335 */
            {8'h00}, /* 0x6334 */
            {8'h00}, /* 0x6333 */
            {8'h00}, /* 0x6332 */
            {8'h00}, /* 0x6331 */
            {8'h00}, /* 0x6330 */
            {8'h00}, /* 0x632f */
            {8'h00}, /* 0x632e */
            {8'h00}, /* 0x632d */
            {8'h00}, /* 0x632c */
            {8'h00}, /* 0x632b */
            {8'h00}, /* 0x632a */
            {8'h00}, /* 0x6329 */
            {8'h00}, /* 0x6328 */
            {8'h00}, /* 0x6327 */
            {8'h00}, /* 0x6326 */
            {8'h00}, /* 0x6325 */
            {8'h00}, /* 0x6324 */
            {8'h00}, /* 0x6323 */
            {8'h00}, /* 0x6322 */
            {8'h00}, /* 0x6321 */
            {8'h00}, /* 0x6320 */
            {8'h00}, /* 0x631f */
            {8'h00}, /* 0x631e */
            {8'h00}, /* 0x631d */
            {8'h00}, /* 0x631c */
            {8'h00}, /* 0x631b */
            {8'h00}, /* 0x631a */
            {8'h00}, /* 0x6319 */
            {8'h00}, /* 0x6318 */
            {8'h00}, /* 0x6317 */
            {8'h00}, /* 0x6316 */
            {8'h00}, /* 0x6315 */
            {8'h00}, /* 0x6314 */
            {8'h00}, /* 0x6313 */
            {8'h00}, /* 0x6312 */
            {8'h00}, /* 0x6311 */
            {8'h00}, /* 0x6310 */
            {8'h00}, /* 0x630f */
            {8'h00}, /* 0x630e */
            {8'h00}, /* 0x630d */
            {8'h00}, /* 0x630c */
            {8'h00}, /* 0x630b */
            {8'h00}, /* 0x630a */
            {8'h00}, /* 0x6309 */
            {8'h00}, /* 0x6308 */
            {8'h00}, /* 0x6307 */
            {8'h00}, /* 0x6306 */
            {8'h00}, /* 0x6305 */
            {8'h00}, /* 0x6304 */
            {8'h00}, /* 0x6303 */
            {8'h00}, /* 0x6302 */
            {8'h00}, /* 0x6301 */
            {8'h00}, /* 0x6300 */
            {8'h00}, /* 0x62ff */
            {8'h00}, /* 0x62fe */
            {8'h00}, /* 0x62fd */
            {8'h00}, /* 0x62fc */
            {8'h00}, /* 0x62fb */
            {8'h00}, /* 0x62fa */
            {8'h00}, /* 0x62f9 */
            {8'h00}, /* 0x62f8 */
            {8'h00}, /* 0x62f7 */
            {8'h00}, /* 0x62f6 */
            {8'h00}, /* 0x62f5 */
            {8'h00}, /* 0x62f4 */
            {8'h00}, /* 0x62f3 */
            {8'h00}, /* 0x62f2 */
            {8'h00}, /* 0x62f1 */
            {8'h00}, /* 0x62f0 */
            {8'h00}, /* 0x62ef */
            {8'h00}, /* 0x62ee */
            {8'h00}, /* 0x62ed */
            {8'h00}, /* 0x62ec */
            {8'h00}, /* 0x62eb */
            {8'h00}, /* 0x62ea */
            {8'h00}, /* 0x62e9 */
            {8'h00}, /* 0x62e8 */
            {8'h00}, /* 0x62e7 */
            {8'h00}, /* 0x62e6 */
            {8'h00}, /* 0x62e5 */
            {8'h00}, /* 0x62e4 */
            {8'h00}, /* 0x62e3 */
            {8'h00}, /* 0x62e2 */
            {8'h00}, /* 0x62e1 */
            {8'h00}, /* 0x62e0 */
            {8'h00}, /* 0x62df */
            {8'h00}, /* 0x62de */
            {8'h00}, /* 0x62dd */
            {8'h00}, /* 0x62dc */
            {8'h00}, /* 0x62db */
            {8'h00}, /* 0x62da */
            {8'h00}, /* 0x62d9 */
            {8'h00}, /* 0x62d8 */
            {8'h00}, /* 0x62d7 */
            {8'h00}, /* 0x62d6 */
            {8'h00}, /* 0x62d5 */
            {8'h00}, /* 0x62d4 */
            {8'h00}, /* 0x62d3 */
            {8'h00}, /* 0x62d2 */
            {8'h00}, /* 0x62d1 */
            {8'h00}, /* 0x62d0 */
            {8'h00}, /* 0x62cf */
            {8'h00}, /* 0x62ce */
            {8'h00}, /* 0x62cd */
            {8'h00}, /* 0x62cc */
            {8'h00}, /* 0x62cb */
            {8'h00}, /* 0x62ca */
            {8'h00}, /* 0x62c9 */
            {8'h00}, /* 0x62c8 */
            {8'h00}, /* 0x62c7 */
            {8'h00}, /* 0x62c6 */
            {8'h00}, /* 0x62c5 */
            {8'h00}, /* 0x62c4 */
            {8'h00}, /* 0x62c3 */
            {8'h00}, /* 0x62c2 */
            {8'h00}, /* 0x62c1 */
            {8'h00}, /* 0x62c0 */
            {8'h00}, /* 0x62bf */
            {8'h00}, /* 0x62be */
            {8'h00}, /* 0x62bd */
            {8'h00}, /* 0x62bc */
            {8'h00}, /* 0x62bb */
            {8'h00}, /* 0x62ba */
            {8'h00}, /* 0x62b9 */
            {8'h00}, /* 0x62b8 */
            {8'h00}, /* 0x62b7 */
            {8'h00}, /* 0x62b6 */
            {8'h00}, /* 0x62b5 */
            {8'h00}, /* 0x62b4 */
            {8'h00}, /* 0x62b3 */
            {8'h00}, /* 0x62b2 */
            {8'h00}, /* 0x62b1 */
            {8'h00}, /* 0x62b0 */
            {8'h00}, /* 0x62af */
            {8'h00}, /* 0x62ae */
            {8'h00}, /* 0x62ad */
            {8'h00}, /* 0x62ac */
            {8'h00}, /* 0x62ab */
            {8'h00}, /* 0x62aa */
            {8'h00}, /* 0x62a9 */
            {8'h00}, /* 0x62a8 */
            {8'h00}, /* 0x62a7 */
            {8'h00}, /* 0x62a6 */
            {8'h00}, /* 0x62a5 */
            {8'h00}, /* 0x62a4 */
            {8'h00}, /* 0x62a3 */
            {8'h00}, /* 0x62a2 */
            {8'h00}, /* 0x62a1 */
            {8'h00}, /* 0x62a0 */
            {8'h00}, /* 0x629f */
            {8'h00}, /* 0x629e */
            {8'h00}, /* 0x629d */
            {8'h00}, /* 0x629c */
            {8'h00}, /* 0x629b */
            {8'h00}, /* 0x629a */
            {8'h00}, /* 0x6299 */
            {8'h00}, /* 0x6298 */
            {8'h00}, /* 0x6297 */
            {8'h00}, /* 0x6296 */
            {8'h00}, /* 0x6295 */
            {8'h00}, /* 0x6294 */
            {8'h00}, /* 0x6293 */
            {8'h00}, /* 0x6292 */
            {8'h00}, /* 0x6291 */
            {8'h00}, /* 0x6290 */
            {8'h00}, /* 0x628f */
            {8'h00}, /* 0x628e */
            {8'h00}, /* 0x628d */
            {8'h00}, /* 0x628c */
            {8'h00}, /* 0x628b */
            {8'h00}, /* 0x628a */
            {8'h00}, /* 0x6289 */
            {8'h00}, /* 0x6288 */
            {8'h00}, /* 0x6287 */
            {8'h00}, /* 0x6286 */
            {8'h00}, /* 0x6285 */
            {8'h00}, /* 0x6284 */
            {8'h00}, /* 0x6283 */
            {8'h00}, /* 0x6282 */
            {8'h00}, /* 0x6281 */
            {8'h00}, /* 0x6280 */
            {8'h00}, /* 0x627f */
            {8'h00}, /* 0x627e */
            {8'h00}, /* 0x627d */
            {8'h00}, /* 0x627c */
            {8'h00}, /* 0x627b */
            {8'h00}, /* 0x627a */
            {8'h00}, /* 0x6279 */
            {8'h00}, /* 0x6278 */
            {8'h00}, /* 0x6277 */
            {8'h00}, /* 0x6276 */
            {8'h00}, /* 0x6275 */
            {8'h00}, /* 0x6274 */
            {8'h00}, /* 0x6273 */
            {8'h00}, /* 0x6272 */
            {8'h00}, /* 0x6271 */
            {8'h00}, /* 0x6270 */
            {8'h00}, /* 0x626f */
            {8'h00}, /* 0x626e */
            {8'h00}, /* 0x626d */
            {8'h00}, /* 0x626c */
            {8'h00}, /* 0x626b */
            {8'h00}, /* 0x626a */
            {8'h00}, /* 0x6269 */
            {8'h00}, /* 0x6268 */
            {8'h00}, /* 0x6267 */
            {8'h00}, /* 0x6266 */
            {8'h00}, /* 0x6265 */
            {8'h00}, /* 0x6264 */
            {8'h00}, /* 0x6263 */
            {8'h00}, /* 0x6262 */
            {8'h00}, /* 0x6261 */
            {8'h00}, /* 0x6260 */
            {8'h00}, /* 0x625f */
            {8'h00}, /* 0x625e */
            {8'h00}, /* 0x625d */
            {8'h00}, /* 0x625c */
            {8'h00}, /* 0x625b */
            {8'h00}, /* 0x625a */
            {8'h00}, /* 0x6259 */
            {8'h00}, /* 0x6258 */
            {8'h00}, /* 0x6257 */
            {8'h00}, /* 0x6256 */
            {8'h00}, /* 0x6255 */
            {8'h00}, /* 0x6254 */
            {8'h00}, /* 0x6253 */
            {8'h00}, /* 0x6252 */
            {8'h00}, /* 0x6251 */
            {8'h00}, /* 0x6250 */
            {8'h00}, /* 0x624f */
            {8'h00}, /* 0x624e */
            {8'h00}, /* 0x624d */
            {8'h00}, /* 0x624c */
            {8'h00}, /* 0x624b */
            {8'h00}, /* 0x624a */
            {8'h00}, /* 0x6249 */
            {8'h00}, /* 0x6248 */
            {8'h00}, /* 0x6247 */
            {8'h00}, /* 0x6246 */
            {8'h00}, /* 0x6245 */
            {8'h00}, /* 0x6244 */
            {8'h00}, /* 0x6243 */
            {8'h00}, /* 0x6242 */
            {8'h00}, /* 0x6241 */
            {8'h00}, /* 0x6240 */
            {8'h00}, /* 0x623f */
            {8'h00}, /* 0x623e */
            {8'h00}, /* 0x623d */
            {8'h00}, /* 0x623c */
            {8'h00}, /* 0x623b */
            {8'h00}, /* 0x623a */
            {8'h00}, /* 0x6239 */
            {8'h00}, /* 0x6238 */
            {8'h00}, /* 0x6237 */
            {8'h00}, /* 0x6236 */
            {8'h00}, /* 0x6235 */
            {8'h00}, /* 0x6234 */
            {8'h00}, /* 0x6233 */
            {8'h00}, /* 0x6232 */
            {8'h00}, /* 0x6231 */
            {8'h00}, /* 0x6230 */
            {8'h00}, /* 0x622f */
            {8'h00}, /* 0x622e */
            {8'h00}, /* 0x622d */
            {8'h00}, /* 0x622c */
            {8'h00}, /* 0x622b */
            {8'h00}, /* 0x622a */
            {8'h00}, /* 0x6229 */
            {8'h00}, /* 0x6228 */
            {8'h00}, /* 0x6227 */
            {8'h00}, /* 0x6226 */
            {8'h00}, /* 0x6225 */
            {8'h00}, /* 0x6224 */
            {8'h00}, /* 0x6223 */
            {8'h00}, /* 0x6222 */
            {8'h00}, /* 0x6221 */
            {8'h00}, /* 0x6220 */
            {8'h00}, /* 0x621f */
            {8'h00}, /* 0x621e */
            {8'h00}, /* 0x621d */
            {8'h00}, /* 0x621c */
            {8'h00}, /* 0x621b */
            {8'h00}, /* 0x621a */
            {8'h00}, /* 0x6219 */
            {8'h00}, /* 0x6218 */
            {8'h00}, /* 0x6217 */
            {8'h00}, /* 0x6216 */
            {8'h00}, /* 0x6215 */
            {8'h00}, /* 0x6214 */
            {8'h00}, /* 0x6213 */
            {8'h00}, /* 0x6212 */
            {8'h00}, /* 0x6211 */
            {8'h00}, /* 0x6210 */
            {8'h00}, /* 0x620f */
            {8'h00}, /* 0x620e */
            {8'h00}, /* 0x620d */
            {8'h00}, /* 0x620c */
            {8'h00}, /* 0x620b */
            {8'h00}, /* 0x620a */
            {8'h00}, /* 0x6209 */
            {8'h00}, /* 0x6208 */
            {8'h00}, /* 0x6207 */
            {8'h00}, /* 0x6206 */
            {8'h00}, /* 0x6205 */
            {8'h00}, /* 0x6204 */
            {8'h00}, /* 0x6203 */
            {8'h00}, /* 0x6202 */
            {8'h00}, /* 0x6201 */
            {8'h00}, /* 0x6200 */
            {8'h00}, /* 0x61ff */
            {8'h00}, /* 0x61fe */
            {8'h00}, /* 0x61fd */
            {8'h00}, /* 0x61fc */
            {8'h00}, /* 0x61fb */
            {8'h00}, /* 0x61fa */
            {8'h00}, /* 0x61f9 */
            {8'h00}, /* 0x61f8 */
            {8'h00}, /* 0x61f7 */
            {8'h00}, /* 0x61f6 */
            {8'h00}, /* 0x61f5 */
            {8'h00}, /* 0x61f4 */
            {8'h00}, /* 0x61f3 */
            {8'h00}, /* 0x61f2 */
            {8'h00}, /* 0x61f1 */
            {8'h00}, /* 0x61f0 */
            {8'h00}, /* 0x61ef */
            {8'h00}, /* 0x61ee */
            {8'h00}, /* 0x61ed */
            {8'h00}, /* 0x61ec */
            {8'h00}, /* 0x61eb */
            {8'h00}, /* 0x61ea */
            {8'h00}, /* 0x61e9 */
            {8'h00}, /* 0x61e8 */
            {8'h00}, /* 0x61e7 */
            {8'h00}, /* 0x61e6 */
            {8'h00}, /* 0x61e5 */
            {8'h00}, /* 0x61e4 */
            {8'h00}, /* 0x61e3 */
            {8'h00}, /* 0x61e2 */
            {8'h00}, /* 0x61e1 */
            {8'h00}, /* 0x61e0 */
            {8'h00}, /* 0x61df */
            {8'h00}, /* 0x61de */
            {8'h00}, /* 0x61dd */
            {8'h00}, /* 0x61dc */
            {8'h00}, /* 0x61db */
            {8'h00}, /* 0x61da */
            {8'h00}, /* 0x61d9 */
            {8'h00}, /* 0x61d8 */
            {8'h00}, /* 0x61d7 */
            {8'h00}, /* 0x61d6 */
            {8'h00}, /* 0x61d5 */
            {8'h00}, /* 0x61d4 */
            {8'h00}, /* 0x61d3 */
            {8'h00}, /* 0x61d2 */
            {8'h00}, /* 0x61d1 */
            {8'h00}, /* 0x61d0 */
            {8'h00}, /* 0x61cf */
            {8'h00}, /* 0x61ce */
            {8'h00}, /* 0x61cd */
            {8'h00}, /* 0x61cc */
            {8'h00}, /* 0x61cb */
            {8'h00}, /* 0x61ca */
            {8'h00}, /* 0x61c9 */
            {8'h00}, /* 0x61c8 */
            {8'h00}, /* 0x61c7 */
            {8'h00}, /* 0x61c6 */
            {8'h00}, /* 0x61c5 */
            {8'h00}, /* 0x61c4 */
            {8'h00}, /* 0x61c3 */
            {8'h00}, /* 0x61c2 */
            {8'h00}, /* 0x61c1 */
            {8'h00}, /* 0x61c0 */
            {8'h00}, /* 0x61bf */
            {8'h00}, /* 0x61be */
            {8'h00}, /* 0x61bd */
            {8'h00}, /* 0x61bc */
            {8'h00}, /* 0x61bb */
            {8'h00}, /* 0x61ba */
            {8'h00}, /* 0x61b9 */
            {8'h00}, /* 0x61b8 */
            {8'h00}, /* 0x61b7 */
            {8'h00}, /* 0x61b6 */
            {8'h00}, /* 0x61b5 */
            {8'h00}, /* 0x61b4 */
            {8'h00}, /* 0x61b3 */
            {8'h00}, /* 0x61b2 */
            {8'h00}, /* 0x61b1 */
            {8'h00}, /* 0x61b0 */
            {8'h00}, /* 0x61af */
            {8'h00}, /* 0x61ae */
            {8'h00}, /* 0x61ad */
            {8'h00}, /* 0x61ac */
            {8'h00}, /* 0x61ab */
            {8'h00}, /* 0x61aa */
            {8'h00}, /* 0x61a9 */
            {8'h00}, /* 0x61a8 */
            {8'h00}, /* 0x61a7 */
            {8'h00}, /* 0x61a6 */
            {8'h00}, /* 0x61a5 */
            {8'h00}, /* 0x61a4 */
            {8'h00}, /* 0x61a3 */
            {8'h00}, /* 0x61a2 */
            {8'h00}, /* 0x61a1 */
            {8'h00}, /* 0x61a0 */
            {8'h00}, /* 0x619f */
            {8'h00}, /* 0x619e */
            {8'h00}, /* 0x619d */
            {8'h00}, /* 0x619c */
            {8'h00}, /* 0x619b */
            {8'h00}, /* 0x619a */
            {8'h00}, /* 0x6199 */
            {8'h00}, /* 0x6198 */
            {8'h00}, /* 0x6197 */
            {8'h00}, /* 0x6196 */
            {8'h00}, /* 0x6195 */
            {8'h00}, /* 0x6194 */
            {8'h00}, /* 0x6193 */
            {8'h00}, /* 0x6192 */
            {8'h00}, /* 0x6191 */
            {8'h00}, /* 0x6190 */
            {8'h00}, /* 0x618f */
            {8'h00}, /* 0x618e */
            {8'h00}, /* 0x618d */
            {8'h00}, /* 0x618c */
            {8'h00}, /* 0x618b */
            {8'h00}, /* 0x618a */
            {8'h00}, /* 0x6189 */
            {8'h00}, /* 0x6188 */
            {8'h00}, /* 0x6187 */
            {8'h00}, /* 0x6186 */
            {8'h00}, /* 0x6185 */
            {8'h00}, /* 0x6184 */
            {8'h00}, /* 0x6183 */
            {8'h00}, /* 0x6182 */
            {8'h00}, /* 0x6181 */
            {8'h00}, /* 0x6180 */
            {8'h00}, /* 0x617f */
            {8'h00}, /* 0x617e */
            {8'h00}, /* 0x617d */
            {8'h00}, /* 0x617c */
            {8'h00}, /* 0x617b */
            {8'h00}, /* 0x617a */
            {8'h00}, /* 0x6179 */
            {8'h00}, /* 0x6178 */
            {8'h00}, /* 0x6177 */
            {8'h00}, /* 0x6176 */
            {8'h00}, /* 0x6175 */
            {8'h00}, /* 0x6174 */
            {8'h00}, /* 0x6173 */
            {8'h00}, /* 0x6172 */
            {8'h00}, /* 0x6171 */
            {8'h00}, /* 0x6170 */
            {8'h00}, /* 0x616f */
            {8'h00}, /* 0x616e */
            {8'h00}, /* 0x616d */
            {8'h00}, /* 0x616c */
            {8'h00}, /* 0x616b */
            {8'h00}, /* 0x616a */
            {8'h00}, /* 0x6169 */
            {8'h00}, /* 0x6168 */
            {8'h00}, /* 0x6167 */
            {8'h00}, /* 0x6166 */
            {8'h00}, /* 0x6165 */
            {8'h00}, /* 0x6164 */
            {8'h00}, /* 0x6163 */
            {8'h00}, /* 0x6162 */
            {8'h00}, /* 0x6161 */
            {8'h00}, /* 0x6160 */
            {8'h00}, /* 0x615f */
            {8'h00}, /* 0x615e */
            {8'h00}, /* 0x615d */
            {8'h00}, /* 0x615c */
            {8'h00}, /* 0x615b */
            {8'h00}, /* 0x615a */
            {8'h00}, /* 0x6159 */
            {8'h00}, /* 0x6158 */
            {8'h00}, /* 0x6157 */
            {8'h00}, /* 0x6156 */
            {8'h00}, /* 0x6155 */
            {8'h00}, /* 0x6154 */
            {8'h00}, /* 0x6153 */
            {8'h00}, /* 0x6152 */
            {8'h00}, /* 0x6151 */
            {8'h00}, /* 0x6150 */
            {8'h00}, /* 0x614f */
            {8'h00}, /* 0x614e */
            {8'h00}, /* 0x614d */
            {8'h00}, /* 0x614c */
            {8'h00}, /* 0x614b */
            {8'h00}, /* 0x614a */
            {8'h00}, /* 0x6149 */
            {8'h00}, /* 0x6148 */
            {8'h00}, /* 0x6147 */
            {8'h00}, /* 0x6146 */
            {8'h00}, /* 0x6145 */
            {8'h00}, /* 0x6144 */
            {8'h00}, /* 0x6143 */
            {8'h00}, /* 0x6142 */
            {8'h00}, /* 0x6141 */
            {8'h00}, /* 0x6140 */
            {8'h00}, /* 0x613f */
            {8'h00}, /* 0x613e */
            {8'h00}, /* 0x613d */
            {8'h00}, /* 0x613c */
            {8'h00}, /* 0x613b */
            {8'h00}, /* 0x613a */
            {8'h00}, /* 0x6139 */
            {8'h00}, /* 0x6138 */
            {8'h00}, /* 0x6137 */
            {8'h00}, /* 0x6136 */
            {8'h00}, /* 0x6135 */
            {8'h00}, /* 0x6134 */
            {8'h00}, /* 0x6133 */
            {8'h00}, /* 0x6132 */
            {8'h00}, /* 0x6131 */
            {8'h00}, /* 0x6130 */
            {8'h00}, /* 0x612f */
            {8'h00}, /* 0x612e */
            {8'h00}, /* 0x612d */
            {8'h00}, /* 0x612c */
            {8'h00}, /* 0x612b */
            {8'h00}, /* 0x612a */
            {8'h00}, /* 0x6129 */
            {8'h00}, /* 0x6128 */
            {8'h00}, /* 0x6127 */
            {8'h00}, /* 0x6126 */
            {8'h00}, /* 0x6125 */
            {8'h00}, /* 0x6124 */
            {8'h00}, /* 0x6123 */
            {8'h00}, /* 0x6122 */
            {8'h00}, /* 0x6121 */
            {8'h00}, /* 0x6120 */
            {8'h00}, /* 0x611f */
            {8'h00}, /* 0x611e */
            {8'h00}, /* 0x611d */
            {8'h00}, /* 0x611c */
            {8'h00}, /* 0x611b */
            {8'h00}, /* 0x611a */
            {8'h00}, /* 0x6119 */
            {8'h00}, /* 0x6118 */
            {8'h00}, /* 0x6117 */
            {8'h00}, /* 0x6116 */
            {8'h00}, /* 0x6115 */
            {8'h00}, /* 0x6114 */
            {8'h00}, /* 0x6113 */
            {8'h00}, /* 0x6112 */
            {8'h00}, /* 0x6111 */
            {8'h00}, /* 0x6110 */
            {8'h00}, /* 0x610f */
            {8'h00}, /* 0x610e */
            {8'h00}, /* 0x610d */
            {8'h00}, /* 0x610c */
            {8'h00}, /* 0x610b */
            {8'h00}, /* 0x610a */
            {8'h00}, /* 0x6109 */
            {8'h00}, /* 0x6108 */
            {8'h00}, /* 0x6107 */
            {8'h00}, /* 0x6106 */
            {8'h00}, /* 0x6105 */
            {8'h00}, /* 0x6104 */
            {8'h00}, /* 0x6103 */
            {8'h00}, /* 0x6102 */
            {8'h00}, /* 0x6101 */
            {8'h00}, /* 0x6100 */
            {8'h00}, /* 0x60ff */
            {8'h00}, /* 0x60fe */
            {8'h00}, /* 0x60fd */
            {8'h00}, /* 0x60fc */
            {8'h00}, /* 0x60fb */
            {8'h00}, /* 0x60fa */
            {8'h00}, /* 0x60f9 */
            {8'h00}, /* 0x60f8 */
            {8'h00}, /* 0x60f7 */
            {8'h00}, /* 0x60f6 */
            {8'h00}, /* 0x60f5 */
            {8'h00}, /* 0x60f4 */
            {8'h00}, /* 0x60f3 */
            {8'h00}, /* 0x60f2 */
            {8'h00}, /* 0x60f1 */
            {8'h00}, /* 0x60f0 */
            {8'h00}, /* 0x60ef */
            {8'h00}, /* 0x60ee */
            {8'h00}, /* 0x60ed */
            {8'h00}, /* 0x60ec */
            {8'h00}, /* 0x60eb */
            {8'h00}, /* 0x60ea */
            {8'h00}, /* 0x60e9 */
            {8'h00}, /* 0x60e8 */
            {8'h00}, /* 0x60e7 */
            {8'h00}, /* 0x60e6 */
            {8'h00}, /* 0x60e5 */
            {8'h00}, /* 0x60e4 */
            {8'h00}, /* 0x60e3 */
            {8'h00}, /* 0x60e2 */
            {8'h00}, /* 0x60e1 */
            {8'h00}, /* 0x60e0 */
            {8'h00}, /* 0x60df */
            {8'h00}, /* 0x60de */
            {8'h00}, /* 0x60dd */
            {8'h00}, /* 0x60dc */
            {8'h00}, /* 0x60db */
            {8'h00}, /* 0x60da */
            {8'h00}, /* 0x60d9 */
            {8'h00}, /* 0x60d8 */
            {8'h00}, /* 0x60d7 */
            {8'h00}, /* 0x60d6 */
            {8'h00}, /* 0x60d5 */
            {8'h00}, /* 0x60d4 */
            {8'h00}, /* 0x60d3 */
            {8'h00}, /* 0x60d2 */
            {8'h00}, /* 0x60d1 */
            {8'h00}, /* 0x60d0 */
            {8'h00}, /* 0x60cf */
            {8'h00}, /* 0x60ce */
            {8'h00}, /* 0x60cd */
            {8'h00}, /* 0x60cc */
            {8'h00}, /* 0x60cb */
            {8'h00}, /* 0x60ca */
            {8'h00}, /* 0x60c9 */
            {8'h00}, /* 0x60c8 */
            {8'h00}, /* 0x60c7 */
            {8'h00}, /* 0x60c6 */
            {8'h00}, /* 0x60c5 */
            {8'h00}, /* 0x60c4 */
            {8'h00}, /* 0x60c3 */
            {8'h00}, /* 0x60c2 */
            {8'h00}, /* 0x60c1 */
            {8'h00}, /* 0x60c0 */
            {8'h00}, /* 0x60bf */
            {8'h00}, /* 0x60be */
            {8'h00}, /* 0x60bd */
            {8'h00}, /* 0x60bc */
            {8'h00}, /* 0x60bb */
            {8'h00}, /* 0x60ba */
            {8'h00}, /* 0x60b9 */
            {8'h00}, /* 0x60b8 */
            {8'h00}, /* 0x60b7 */
            {8'h00}, /* 0x60b6 */
            {8'h00}, /* 0x60b5 */
            {8'h00}, /* 0x60b4 */
            {8'h00}, /* 0x60b3 */
            {8'h00}, /* 0x60b2 */
            {8'h00}, /* 0x60b1 */
            {8'h00}, /* 0x60b0 */
            {8'h00}, /* 0x60af */
            {8'h00}, /* 0x60ae */
            {8'h00}, /* 0x60ad */
            {8'h00}, /* 0x60ac */
            {8'h00}, /* 0x60ab */
            {8'h00}, /* 0x60aa */
            {8'h00}, /* 0x60a9 */
            {8'h00}, /* 0x60a8 */
            {8'h00}, /* 0x60a7 */
            {8'h00}, /* 0x60a6 */
            {8'h00}, /* 0x60a5 */
            {8'h00}, /* 0x60a4 */
            {8'h00}, /* 0x60a3 */
            {8'h00}, /* 0x60a2 */
            {8'h00}, /* 0x60a1 */
            {8'h00}, /* 0x60a0 */
            {8'h00}, /* 0x609f */
            {8'h00}, /* 0x609e */
            {8'h00}, /* 0x609d */
            {8'h00}, /* 0x609c */
            {8'h00}, /* 0x609b */
            {8'h00}, /* 0x609a */
            {8'h00}, /* 0x6099 */
            {8'h00}, /* 0x6098 */
            {8'h00}, /* 0x6097 */
            {8'h00}, /* 0x6096 */
            {8'h00}, /* 0x6095 */
            {8'h00}, /* 0x6094 */
            {8'h00}, /* 0x6093 */
            {8'h00}, /* 0x6092 */
            {8'h00}, /* 0x6091 */
            {8'h00}, /* 0x6090 */
            {8'h00}, /* 0x608f */
            {8'h00}, /* 0x608e */
            {8'h00}, /* 0x608d */
            {8'h00}, /* 0x608c */
            {8'h00}, /* 0x608b */
            {8'h00}, /* 0x608a */
            {8'h00}, /* 0x6089 */
            {8'h00}, /* 0x6088 */
            {8'h00}, /* 0x6087 */
            {8'h00}, /* 0x6086 */
            {8'h00}, /* 0x6085 */
            {8'h00}, /* 0x6084 */
            {8'h00}, /* 0x6083 */
            {8'h00}, /* 0x6082 */
            {8'h00}, /* 0x6081 */
            {8'h00}, /* 0x6080 */
            {8'h00}, /* 0x607f */
            {8'h00}, /* 0x607e */
            {8'h00}, /* 0x607d */
            {8'h00}, /* 0x607c */
            {8'h00}, /* 0x607b */
            {8'h00}, /* 0x607a */
            {8'h00}, /* 0x6079 */
            {8'h00}, /* 0x6078 */
            {8'h00}, /* 0x6077 */
            {8'h00}, /* 0x6076 */
            {8'h00}, /* 0x6075 */
            {8'h00}, /* 0x6074 */
            {8'h00}, /* 0x6073 */
            {8'h00}, /* 0x6072 */
            {8'h00}, /* 0x6071 */
            {8'h00}, /* 0x6070 */
            {8'h00}, /* 0x606f */
            {8'h00}, /* 0x606e */
            {8'h00}, /* 0x606d */
            {8'h00}, /* 0x606c */
            {8'h00}, /* 0x606b */
            {8'h00}, /* 0x606a */
            {8'h00}, /* 0x6069 */
            {8'h00}, /* 0x6068 */
            {8'h00}, /* 0x6067 */
            {8'h00}, /* 0x6066 */
            {8'h00}, /* 0x6065 */
            {8'h00}, /* 0x6064 */
            {8'h00}, /* 0x6063 */
            {8'h00}, /* 0x6062 */
            {8'h00}, /* 0x6061 */
            {8'h00}, /* 0x6060 */
            {8'h00}, /* 0x605f */
            {8'h00}, /* 0x605e */
            {8'h00}, /* 0x605d */
            {8'h00}, /* 0x605c */
            {8'h00}, /* 0x605b */
            {8'h00}, /* 0x605a */
            {8'h00}, /* 0x6059 */
            {8'h00}, /* 0x6058 */
            {8'h00}, /* 0x6057 */
            {8'h00}, /* 0x6056 */
            {8'h00}, /* 0x6055 */
            {8'h00}, /* 0x6054 */
            {8'h00}, /* 0x6053 */
            {8'h00}, /* 0x6052 */
            {8'h00}, /* 0x6051 */
            {8'h00}, /* 0x6050 */
            {8'h00}, /* 0x604f */
            {8'h00}, /* 0x604e */
            {8'h00}, /* 0x604d */
            {8'h00}, /* 0x604c */
            {8'h00}, /* 0x604b */
            {8'h00}, /* 0x604a */
            {8'h00}, /* 0x6049 */
            {8'h00}, /* 0x6048 */
            {8'h00}, /* 0x6047 */
            {8'h00}, /* 0x6046 */
            {8'h00}, /* 0x6045 */
            {8'h00}, /* 0x6044 */
            {8'h00}, /* 0x6043 */
            {8'h00}, /* 0x6042 */
            {8'h00}, /* 0x6041 */
            {8'h00}, /* 0x6040 */
            {8'h00}, /* 0x603f */
            {8'h00}, /* 0x603e */
            {8'h00}, /* 0x603d */
            {8'h00}, /* 0x603c */
            {8'h00}, /* 0x603b */
            {8'h00}, /* 0x603a */
            {8'h00}, /* 0x6039 */
            {8'h00}, /* 0x6038 */
            {8'h00}, /* 0x6037 */
            {8'h00}, /* 0x6036 */
            {8'h00}, /* 0x6035 */
            {8'h00}, /* 0x6034 */
            {8'h00}, /* 0x6033 */
            {8'h00}, /* 0x6032 */
            {8'h00}, /* 0x6031 */
            {8'h00}, /* 0x6030 */
            {8'h00}, /* 0x602f */
            {8'h00}, /* 0x602e */
            {8'h00}, /* 0x602d */
            {8'h00}, /* 0x602c */
            {8'h00}, /* 0x602b */
            {8'h00}, /* 0x602a */
            {8'h00}, /* 0x6029 */
            {8'h00}, /* 0x6028 */
            {8'h00}, /* 0x6027 */
            {8'h00}, /* 0x6026 */
            {8'h00}, /* 0x6025 */
            {8'h00}, /* 0x6024 */
            {8'h00}, /* 0x6023 */
            {8'h00}, /* 0x6022 */
            {8'h00}, /* 0x6021 */
            {8'h00}, /* 0x6020 */
            {8'h00}, /* 0x601f */
            {8'h00}, /* 0x601e */
            {8'h00}, /* 0x601d */
            {8'h00}, /* 0x601c */
            {8'h00}, /* 0x601b */
            {8'h00}, /* 0x601a */
            {8'h00}, /* 0x6019 */
            {8'h00}, /* 0x6018 */
            {8'h00}, /* 0x6017 */
            {8'h00}, /* 0x6016 */
            {8'h00}, /* 0x6015 */
            {8'h00}, /* 0x6014 */
            {8'h00}, /* 0x6013 */
            {8'h00}, /* 0x6012 */
            {8'h00}, /* 0x6011 */
            {8'h00}, /* 0x6010 */
            {8'h00}, /* 0x600f */
            {8'h00}, /* 0x600e */
            {8'h00}, /* 0x600d */
            {8'h00}, /* 0x600c */
            {8'h00}, /* 0x600b */
            {8'h00}, /* 0x600a */
            {8'h00}, /* 0x6009 */
            {8'h00}, /* 0x6008 */
            {8'h00}, /* 0x6007 */
            {8'h00}, /* 0x6006 */
            {8'h00}, /* 0x6005 */
            {8'h00}, /* 0x6004 */
            {8'h00}, /* 0x6003 */
            {8'h00}, /* 0x6002 */
            {8'h00}, /* 0x6001 */
            {8'h00}, /* 0x6000 */
            {8'h00}, /* 0x5fff */
            {8'h00}, /* 0x5ffe */
            {8'h00}, /* 0x5ffd */
            {8'h00}, /* 0x5ffc */
            {8'h00}, /* 0x5ffb */
            {8'h00}, /* 0x5ffa */
            {8'h00}, /* 0x5ff9 */
            {8'h00}, /* 0x5ff8 */
            {8'h00}, /* 0x5ff7 */
            {8'h00}, /* 0x5ff6 */
            {8'h00}, /* 0x5ff5 */
            {8'h00}, /* 0x5ff4 */
            {8'h00}, /* 0x5ff3 */
            {8'h00}, /* 0x5ff2 */
            {8'h00}, /* 0x5ff1 */
            {8'h00}, /* 0x5ff0 */
            {8'h00}, /* 0x5fef */
            {8'h00}, /* 0x5fee */
            {8'h00}, /* 0x5fed */
            {8'h00}, /* 0x5fec */
            {8'h00}, /* 0x5feb */
            {8'h00}, /* 0x5fea */
            {8'h00}, /* 0x5fe9 */
            {8'h00}, /* 0x5fe8 */
            {8'h00}, /* 0x5fe7 */
            {8'h00}, /* 0x5fe6 */
            {8'h00}, /* 0x5fe5 */
            {8'h00}, /* 0x5fe4 */
            {8'h00}, /* 0x5fe3 */
            {8'h00}, /* 0x5fe2 */
            {8'h00}, /* 0x5fe1 */
            {8'h00}, /* 0x5fe0 */
            {8'h00}, /* 0x5fdf */
            {8'h00}, /* 0x5fde */
            {8'h00}, /* 0x5fdd */
            {8'h00}, /* 0x5fdc */
            {8'h00}, /* 0x5fdb */
            {8'h00}, /* 0x5fda */
            {8'h00}, /* 0x5fd9 */
            {8'h00}, /* 0x5fd8 */
            {8'h00}, /* 0x5fd7 */
            {8'h00}, /* 0x5fd6 */
            {8'h00}, /* 0x5fd5 */
            {8'h00}, /* 0x5fd4 */
            {8'h00}, /* 0x5fd3 */
            {8'h00}, /* 0x5fd2 */
            {8'h00}, /* 0x5fd1 */
            {8'h00}, /* 0x5fd0 */
            {8'h00}, /* 0x5fcf */
            {8'h00}, /* 0x5fce */
            {8'h00}, /* 0x5fcd */
            {8'h00}, /* 0x5fcc */
            {8'h00}, /* 0x5fcb */
            {8'h00}, /* 0x5fca */
            {8'h00}, /* 0x5fc9 */
            {8'h00}, /* 0x5fc8 */
            {8'h00}, /* 0x5fc7 */
            {8'h00}, /* 0x5fc6 */
            {8'h00}, /* 0x5fc5 */
            {8'h00}, /* 0x5fc4 */
            {8'h00}, /* 0x5fc3 */
            {8'h00}, /* 0x5fc2 */
            {8'h00}, /* 0x5fc1 */
            {8'h00}, /* 0x5fc0 */
            {8'h00}, /* 0x5fbf */
            {8'h00}, /* 0x5fbe */
            {8'h00}, /* 0x5fbd */
            {8'h00}, /* 0x5fbc */
            {8'h00}, /* 0x5fbb */
            {8'h00}, /* 0x5fba */
            {8'h00}, /* 0x5fb9 */
            {8'h00}, /* 0x5fb8 */
            {8'h00}, /* 0x5fb7 */
            {8'h00}, /* 0x5fb6 */
            {8'h00}, /* 0x5fb5 */
            {8'h00}, /* 0x5fb4 */
            {8'h00}, /* 0x5fb3 */
            {8'h00}, /* 0x5fb2 */
            {8'h00}, /* 0x5fb1 */
            {8'h00}, /* 0x5fb0 */
            {8'h00}, /* 0x5faf */
            {8'h00}, /* 0x5fae */
            {8'h00}, /* 0x5fad */
            {8'h00}, /* 0x5fac */
            {8'h00}, /* 0x5fab */
            {8'h00}, /* 0x5faa */
            {8'h00}, /* 0x5fa9 */
            {8'h00}, /* 0x5fa8 */
            {8'h00}, /* 0x5fa7 */
            {8'h00}, /* 0x5fa6 */
            {8'h00}, /* 0x5fa5 */
            {8'h00}, /* 0x5fa4 */
            {8'h00}, /* 0x5fa3 */
            {8'h00}, /* 0x5fa2 */
            {8'h00}, /* 0x5fa1 */
            {8'h00}, /* 0x5fa0 */
            {8'h00}, /* 0x5f9f */
            {8'h00}, /* 0x5f9e */
            {8'h00}, /* 0x5f9d */
            {8'h00}, /* 0x5f9c */
            {8'h00}, /* 0x5f9b */
            {8'h00}, /* 0x5f9a */
            {8'h00}, /* 0x5f99 */
            {8'h00}, /* 0x5f98 */
            {8'h00}, /* 0x5f97 */
            {8'h00}, /* 0x5f96 */
            {8'h00}, /* 0x5f95 */
            {8'h00}, /* 0x5f94 */
            {8'h00}, /* 0x5f93 */
            {8'h00}, /* 0x5f92 */
            {8'h00}, /* 0x5f91 */
            {8'h00}, /* 0x5f90 */
            {8'h00}, /* 0x5f8f */
            {8'h00}, /* 0x5f8e */
            {8'h00}, /* 0x5f8d */
            {8'h00}, /* 0x5f8c */
            {8'h00}, /* 0x5f8b */
            {8'h00}, /* 0x5f8a */
            {8'h00}, /* 0x5f89 */
            {8'h00}, /* 0x5f88 */
            {8'h00}, /* 0x5f87 */
            {8'h00}, /* 0x5f86 */
            {8'h00}, /* 0x5f85 */
            {8'h00}, /* 0x5f84 */
            {8'h00}, /* 0x5f83 */
            {8'h00}, /* 0x5f82 */
            {8'h00}, /* 0x5f81 */
            {8'h00}, /* 0x5f80 */
            {8'h00}, /* 0x5f7f */
            {8'h00}, /* 0x5f7e */
            {8'h00}, /* 0x5f7d */
            {8'h00}, /* 0x5f7c */
            {8'h00}, /* 0x5f7b */
            {8'h00}, /* 0x5f7a */
            {8'h00}, /* 0x5f79 */
            {8'h00}, /* 0x5f78 */
            {8'h00}, /* 0x5f77 */
            {8'h00}, /* 0x5f76 */
            {8'h00}, /* 0x5f75 */
            {8'h00}, /* 0x5f74 */
            {8'h00}, /* 0x5f73 */
            {8'h00}, /* 0x5f72 */
            {8'h00}, /* 0x5f71 */
            {8'h00}, /* 0x5f70 */
            {8'h00}, /* 0x5f6f */
            {8'h00}, /* 0x5f6e */
            {8'h00}, /* 0x5f6d */
            {8'h00}, /* 0x5f6c */
            {8'h00}, /* 0x5f6b */
            {8'h00}, /* 0x5f6a */
            {8'h00}, /* 0x5f69 */
            {8'h00}, /* 0x5f68 */
            {8'h00}, /* 0x5f67 */
            {8'h00}, /* 0x5f66 */
            {8'h00}, /* 0x5f65 */
            {8'h00}, /* 0x5f64 */
            {8'h00}, /* 0x5f63 */
            {8'h00}, /* 0x5f62 */
            {8'h00}, /* 0x5f61 */
            {8'h00}, /* 0x5f60 */
            {8'h00}, /* 0x5f5f */
            {8'h00}, /* 0x5f5e */
            {8'h00}, /* 0x5f5d */
            {8'h00}, /* 0x5f5c */
            {8'h00}, /* 0x5f5b */
            {8'h00}, /* 0x5f5a */
            {8'h00}, /* 0x5f59 */
            {8'h00}, /* 0x5f58 */
            {8'h00}, /* 0x5f57 */
            {8'h00}, /* 0x5f56 */
            {8'h00}, /* 0x5f55 */
            {8'h00}, /* 0x5f54 */
            {8'h00}, /* 0x5f53 */
            {8'h00}, /* 0x5f52 */
            {8'h00}, /* 0x5f51 */
            {8'h00}, /* 0x5f50 */
            {8'h00}, /* 0x5f4f */
            {8'h00}, /* 0x5f4e */
            {8'h00}, /* 0x5f4d */
            {8'h00}, /* 0x5f4c */
            {8'h00}, /* 0x5f4b */
            {8'h00}, /* 0x5f4a */
            {8'h00}, /* 0x5f49 */
            {8'h00}, /* 0x5f48 */
            {8'h00}, /* 0x5f47 */
            {8'h00}, /* 0x5f46 */
            {8'h00}, /* 0x5f45 */
            {8'h00}, /* 0x5f44 */
            {8'h00}, /* 0x5f43 */
            {8'h00}, /* 0x5f42 */
            {8'h00}, /* 0x5f41 */
            {8'h00}, /* 0x5f40 */
            {8'h00}, /* 0x5f3f */
            {8'h00}, /* 0x5f3e */
            {8'h00}, /* 0x5f3d */
            {8'h00}, /* 0x5f3c */
            {8'h00}, /* 0x5f3b */
            {8'h00}, /* 0x5f3a */
            {8'h00}, /* 0x5f39 */
            {8'h00}, /* 0x5f38 */
            {8'h00}, /* 0x5f37 */
            {8'h00}, /* 0x5f36 */
            {8'h00}, /* 0x5f35 */
            {8'h00}, /* 0x5f34 */
            {8'h00}, /* 0x5f33 */
            {8'h00}, /* 0x5f32 */
            {8'h00}, /* 0x5f31 */
            {8'h00}, /* 0x5f30 */
            {8'h00}, /* 0x5f2f */
            {8'h00}, /* 0x5f2e */
            {8'h00}, /* 0x5f2d */
            {8'h00}, /* 0x5f2c */
            {8'h00}, /* 0x5f2b */
            {8'h00}, /* 0x5f2a */
            {8'h00}, /* 0x5f29 */
            {8'h00}, /* 0x5f28 */
            {8'h00}, /* 0x5f27 */
            {8'h00}, /* 0x5f26 */
            {8'h00}, /* 0x5f25 */
            {8'h00}, /* 0x5f24 */
            {8'h00}, /* 0x5f23 */
            {8'h00}, /* 0x5f22 */
            {8'h00}, /* 0x5f21 */
            {8'h00}, /* 0x5f20 */
            {8'h00}, /* 0x5f1f */
            {8'h00}, /* 0x5f1e */
            {8'h00}, /* 0x5f1d */
            {8'h00}, /* 0x5f1c */
            {8'h00}, /* 0x5f1b */
            {8'h00}, /* 0x5f1a */
            {8'h00}, /* 0x5f19 */
            {8'h00}, /* 0x5f18 */
            {8'h00}, /* 0x5f17 */
            {8'h00}, /* 0x5f16 */
            {8'h00}, /* 0x5f15 */
            {8'h00}, /* 0x5f14 */
            {8'h00}, /* 0x5f13 */
            {8'h00}, /* 0x5f12 */
            {8'h00}, /* 0x5f11 */
            {8'h00}, /* 0x5f10 */
            {8'h00}, /* 0x5f0f */
            {8'h00}, /* 0x5f0e */
            {8'h00}, /* 0x5f0d */
            {8'h00}, /* 0x5f0c */
            {8'h00}, /* 0x5f0b */
            {8'h00}, /* 0x5f0a */
            {8'h00}, /* 0x5f09 */
            {8'h00}, /* 0x5f08 */
            {8'h00}, /* 0x5f07 */
            {8'h00}, /* 0x5f06 */
            {8'h00}, /* 0x5f05 */
            {8'h00}, /* 0x5f04 */
            {8'h00}, /* 0x5f03 */
            {8'h00}, /* 0x5f02 */
            {8'h00}, /* 0x5f01 */
            {8'h00}, /* 0x5f00 */
            {8'h00}, /* 0x5eff */
            {8'h00}, /* 0x5efe */
            {8'h00}, /* 0x5efd */
            {8'h00}, /* 0x5efc */
            {8'h00}, /* 0x5efb */
            {8'h00}, /* 0x5efa */
            {8'h00}, /* 0x5ef9 */
            {8'h00}, /* 0x5ef8 */
            {8'h00}, /* 0x5ef7 */
            {8'h00}, /* 0x5ef6 */
            {8'h00}, /* 0x5ef5 */
            {8'h00}, /* 0x5ef4 */
            {8'h00}, /* 0x5ef3 */
            {8'h00}, /* 0x5ef2 */
            {8'h00}, /* 0x5ef1 */
            {8'h00}, /* 0x5ef0 */
            {8'h00}, /* 0x5eef */
            {8'h00}, /* 0x5eee */
            {8'h00}, /* 0x5eed */
            {8'h00}, /* 0x5eec */
            {8'h00}, /* 0x5eeb */
            {8'h00}, /* 0x5eea */
            {8'h00}, /* 0x5ee9 */
            {8'h00}, /* 0x5ee8 */
            {8'h00}, /* 0x5ee7 */
            {8'h00}, /* 0x5ee6 */
            {8'h00}, /* 0x5ee5 */
            {8'h00}, /* 0x5ee4 */
            {8'h00}, /* 0x5ee3 */
            {8'h00}, /* 0x5ee2 */
            {8'h00}, /* 0x5ee1 */
            {8'h00}, /* 0x5ee0 */
            {8'h00}, /* 0x5edf */
            {8'h00}, /* 0x5ede */
            {8'h00}, /* 0x5edd */
            {8'h00}, /* 0x5edc */
            {8'h00}, /* 0x5edb */
            {8'h00}, /* 0x5eda */
            {8'h00}, /* 0x5ed9 */
            {8'h00}, /* 0x5ed8 */
            {8'h00}, /* 0x5ed7 */
            {8'h00}, /* 0x5ed6 */
            {8'h00}, /* 0x5ed5 */
            {8'h00}, /* 0x5ed4 */
            {8'h00}, /* 0x5ed3 */
            {8'h00}, /* 0x5ed2 */
            {8'h00}, /* 0x5ed1 */
            {8'h00}, /* 0x5ed0 */
            {8'h00}, /* 0x5ecf */
            {8'h00}, /* 0x5ece */
            {8'h00}, /* 0x5ecd */
            {8'h00}, /* 0x5ecc */
            {8'h00}, /* 0x5ecb */
            {8'h00}, /* 0x5eca */
            {8'h00}, /* 0x5ec9 */
            {8'h00}, /* 0x5ec8 */
            {8'h00}, /* 0x5ec7 */
            {8'h00}, /* 0x5ec6 */
            {8'h00}, /* 0x5ec5 */
            {8'h00}, /* 0x5ec4 */
            {8'h00}, /* 0x5ec3 */
            {8'h00}, /* 0x5ec2 */
            {8'h00}, /* 0x5ec1 */
            {8'h00}, /* 0x5ec0 */
            {8'h00}, /* 0x5ebf */
            {8'h00}, /* 0x5ebe */
            {8'h00}, /* 0x5ebd */
            {8'h00}, /* 0x5ebc */
            {8'h00}, /* 0x5ebb */
            {8'h00}, /* 0x5eba */
            {8'h00}, /* 0x5eb9 */
            {8'h00}, /* 0x5eb8 */
            {8'h00}, /* 0x5eb7 */
            {8'h00}, /* 0x5eb6 */
            {8'h00}, /* 0x5eb5 */
            {8'h00}, /* 0x5eb4 */
            {8'h00}, /* 0x5eb3 */
            {8'h00}, /* 0x5eb2 */
            {8'h00}, /* 0x5eb1 */
            {8'h00}, /* 0x5eb0 */
            {8'h00}, /* 0x5eaf */
            {8'h00}, /* 0x5eae */
            {8'h00}, /* 0x5ead */
            {8'h00}, /* 0x5eac */
            {8'h00}, /* 0x5eab */
            {8'h00}, /* 0x5eaa */
            {8'h00}, /* 0x5ea9 */
            {8'h00}, /* 0x5ea8 */
            {8'h00}, /* 0x5ea7 */
            {8'h00}, /* 0x5ea6 */
            {8'h00}, /* 0x5ea5 */
            {8'h00}, /* 0x5ea4 */
            {8'h00}, /* 0x5ea3 */
            {8'h00}, /* 0x5ea2 */
            {8'h00}, /* 0x5ea1 */
            {8'h00}, /* 0x5ea0 */
            {8'h00}, /* 0x5e9f */
            {8'h00}, /* 0x5e9e */
            {8'h00}, /* 0x5e9d */
            {8'h00}, /* 0x5e9c */
            {8'h00}, /* 0x5e9b */
            {8'h00}, /* 0x5e9a */
            {8'h00}, /* 0x5e99 */
            {8'h00}, /* 0x5e98 */
            {8'h00}, /* 0x5e97 */
            {8'h00}, /* 0x5e96 */
            {8'h00}, /* 0x5e95 */
            {8'h00}, /* 0x5e94 */
            {8'h00}, /* 0x5e93 */
            {8'h00}, /* 0x5e92 */
            {8'h00}, /* 0x5e91 */
            {8'h00}, /* 0x5e90 */
            {8'h00}, /* 0x5e8f */
            {8'h00}, /* 0x5e8e */
            {8'h00}, /* 0x5e8d */
            {8'h00}, /* 0x5e8c */
            {8'h00}, /* 0x5e8b */
            {8'h00}, /* 0x5e8a */
            {8'h00}, /* 0x5e89 */
            {8'h00}, /* 0x5e88 */
            {8'h00}, /* 0x5e87 */
            {8'h00}, /* 0x5e86 */
            {8'h00}, /* 0x5e85 */
            {8'h00}, /* 0x5e84 */
            {8'h00}, /* 0x5e83 */
            {8'h00}, /* 0x5e82 */
            {8'h00}, /* 0x5e81 */
            {8'h00}, /* 0x5e80 */
            {8'h00}, /* 0x5e7f */
            {8'h00}, /* 0x5e7e */
            {8'h00}, /* 0x5e7d */
            {8'h00}, /* 0x5e7c */
            {8'h00}, /* 0x5e7b */
            {8'h00}, /* 0x5e7a */
            {8'h00}, /* 0x5e79 */
            {8'h00}, /* 0x5e78 */
            {8'h00}, /* 0x5e77 */
            {8'h00}, /* 0x5e76 */
            {8'h00}, /* 0x5e75 */
            {8'h00}, /* 0x5e74 */
            {8'h00}, /* 0x5e73 */
            {8'h00}, /* 0x5e72 */
            {8'h00}, /* 0x5e71 */
            {8'h00}, /* 0x5e70 */
            {8'h00}, /* 0x5e6f */
            {8'h00}, /* 0x5e6e */
            {8'h00}, /* 0x5e6d */
            {8'h00}, /* 0x5e6c */
            {8'h00}, /* 0x5e6b */
            {8'h00}, /* 0x5e6a */
            {8'h00}, /* 0x5e69 */
            {8'h00}, /* 0x5e68 */
            {8'h00}, /* 0x5e67 */
            {8'h00}, /* 0x5e66 */
            {8'h00}, /* 0x5e65 */
            {8'h00}, /* 0x5e64 */
            {8'h00}, /* 0x5e63 */
            {8'h00}, /* 0x5e62 */
            {8'h00}, /* 0x5e61 */
            {8'h00}, /* 0x5e60 */
            {8'h00}, /* 0x5e5f */
            {8'h00}, /* 0x5e5e */
            {8'h00}, /* 0x5e5d */
            {8'h00}, /* 0x5e5c */
            {8'h00}, /* 0x5e5b */
            {8'h00}, /* 0x5e5a */
            {8'h00}, /* 0x5e59 */
            {8'h00}, /* 0x5e58 */
            {8'h00}, /* 0x5e57 */
            {8'h00}, /* 0x5e56 */
            {8'h00}, /* 0x5e55 */
            {8'h00}, /* 0x5e54 */
            {8'h00}, /* 0x5e53 */
            {8'h00}, /* 0x5e52 */
            {8'h00}, /* 0x5e51 */
            {8'h00}, /* 0x5e50 */
            {8'h00}, /* 0x5e4f */
            {8'h00}, /* 0x5e4e */
            {8'h00}, /* 0x5e4d */
            {8'h00}, /* 0x5e4c */
            {8'h00}, /* 0x5e4b */
            {8'h00}, /* 0x5e4a */
            {8'h00}, /* 0x5e49 */
            {8'h00}, /* 0x5e48 */
            {8'h00}, /* 0x5e47 */
            {8'h00}, /* 0x5e46 */
            {8'h00}, /* 0x5e45 */
            {8'h00}, /* 0x5e44 */
            {8'h00}, /* 0x5e43 */
            {8'h00}, /* 0x5e42 */
            {8'h00}, /* 0x5e41 */
            {8'h00}, /* 0x5e40 */
            {8'h00}, /* 0x5e3f */
            {8'h00}, /* 0x5e3e */
            {8'h00}, /* 0x5e3d */
            {8'h00}, /* 0x5e3c */
            {8'h00}, /* 0x5e3b */
            {8'h00}, /* 0x5e3a */
            {8'h00}, /* 0x5e39 */
            {8'h00}, /* 0x5e38 */
            {8'h00}, /* 0x5e37 */
            {8'h00}, /* 0x5e36 */
            {8'h00}, /* 0x5e35 */
            {8'h00}, /* 0x5e34 */
            {8'h00}, /* 0x5e33 */
            {8'h00}, /* 0x5e32 */
            {8'h00}, /* 0x5e31 */
            {8'h00}, /* 0x5e30 */
            {8'h00}, /* 0x5e2f */
            {8'h00}, /* 0x5e2e */
            {8'h00}, /* 0x5e2d */
            {8'h00}, /* 0x5e2c */
            {8'h00}, /* 0x5e2b */
            {8'h00}, /* 0x5e2a */
            {8'h00}, /* 0x5e29 */
            {8'h00}, /* 0x5e28 */
            {8'h00}, /* 0x5e27 */
            {8'h00}, /* 0x5e26 */
            {8'h00}, /* 0x5e25 */
            {8'h00}, /* 0x5e24 */
            {8'h00}, /* 0x5e23 */
            {8'h00}, /* 0x5e22 */
            {8'h00}, /* 0x5e21 */
            {8'h00}, /* 0x5e20 */
            {8'h00}, /* 0x5e1f */
            {8'h00}, /* 0x5e1e */
            {8'h00}, /* 0x5e1d */
            {8'h00}, /* 0x5e1c */
            {8'h00}, /* 0x5e1b */
            {8'h00}, /* 0x5e1a */
            {8'h00}, /* 0x5e19 */
            {8'h00}, /* 0x5e18 */
            {8'h00}, /* 0x5e17 */
            {8'h00}, /* 0x5e16 */
            {8'h00}, /* 0x5e15 */
            {8'h00}, /* 0x5e14 */
            {8'h00}, /* 0x5e13 */
            {8'h00}, /* 0x5e12 */
            {8'h00}, /* 0x5e11 */
            {8'h00}, /* 0x5e10 */
            {8'h00}, /* 0x5e0f */
            {8'h00}, /* 0x5e0e */
            {8'h00}, /* 0x5e0d */
            {8'h00}, /* 0x5e0c */
            {8'h00}, /* 0x5e0b */
            {8'h00}, /* 0x5e0a */
            {8'h00}, /* 0x5e09 */
            {8'h00}, /* 0x5e08 */
            {8'h00}, /* 0x5e07 */
            {8'h00}, /* 0x5e06 */
            {8'h00}, /* 0x5e05 */
            {8'h00}, /* 0x5e04 */
            {8'h00}, /* 0x5e03 */
            {8'h00}, /* 0x5e02 */
            {8'h00}, /* 0x5e01 */
            {8'h00}, /* 0x5e00 */
            {8'h00}, /* 0x5dff */
            {8'h00}, /* 0x5dfe */
            {8'h00}, /* 0x5dfd */
            {8'h00}, /* 0x5dfc */
            {8'h00}, /* 0x5dfb */
            {8'h00}, /* 0x5dfa */
            {8'h00}, /* 0x5df9 */
            {8'h00}, /* 0x5df8 */
            {8'h00}, /* 0x5df7 */
            {8'h00}, /* 0x5df6 */
            {8'h00}, /* 0x5df5 */
            {8'h00}, /* 0x5df4 */
            {8'h00}, /* 0x5df3 */
            {8'h00}, /* 0x5df2 */
            {8'h00}, /* 0x5df1 */
            {8'h00}, /* 0x5df0 */
            {8'h00}, /* 0x5def */
            {8'h00}, /* 0x5dee */
            {8'h00}, /* 0x5ded */
            {8'h00}, /* 0x5dec */
            {8'h00}, /* 0x5deb */
            {8'h00}, /* 0x5dea */
            {8'h00}, /* 0x5de9 */
            {8'h00}, /* 0x5de8 */
            {8'h00}, /* 0x5de7 */
            {8'h00}, /* 0x5de6 */
            {8'h00}, /* 0x5de5 */
            {8'h00}, /* 0x5de4 */
            {8'h00}, /* 0x5de3 */
            {8'h00}, /* 0x5de2 */
            {8'h00}, /* 0x5de1 */
            {8'h00}, /* 0x5de0 */
            {8'h00}, /* 0x5ddf */
            {8'h00}, /* 0x5dde */
            {8'h00}, /* 0x5ddd */
            {8'h00}, /* 0x5ddc */
            {8'h00}, /* 0x5ddb */
            {8'h00}, /* 0x5dda */
            {8'h00}, /* 0x5dd9 */
            {8'h00}, /* 0x5dd8 */
            {8'h00}, /* 0x5dd7 */
            {8'h00}, /* 0x5dd6 */
            {8'h00}, /* 0x5dd5 */
            {8'h00}, /* 0x5dd4 */
            {8'h00}, /* 0x5dd3 */
            {8'h00}, /* 0x5dd2 */
            {8'h00}, /* 0x5dd1 */
            {8'h00}, /* 0x5dd0 */
            {8'h00}, /* 0x5dcf */
            {8'h00}, /* 0x5dce */
            {8'h00}, /* 0x5dcd */
            {8'h00}, /* 0x5dcc */
            {8'h00}, /* 0x5dcb */
            {8'h00}, /* 0x5dca */
            {8'h00}, /* 0x5dc9 */
            {8'h00}, /* 0x5dc8 */
            {8'h00}, /* 0x5dc7 */
            {8'h00}, /* 0x5dc6 */
            {8'h00}, /* 0x5dc5 */
            {8'h00}, /* 0x5dc4 */
            {8'h00}, /* 0x5dc3 */
            {8'h00}, /* 0x5dc2 */
            {8'h00}, /* 0x5dc1 */
            {8'h00}, /* 0x5dc0 */
            {8'h00}, /* 0x5dbf */
            {8'h00}, /* 0x5dbe */
            {8'h00}, /* 0x5dbd */
            {8'h00}, /* 0x5dbc */
            {8'h00}, /* 0x5dbb */
            {8'h00}, /* 0x5dba */
            {8'h00}, /* 0x5db9 */
            {8'h00}, /* 0x5db8 */
            {8'h00}, /* 0x5db7 */
            {8'h00}, /* 0x5db6 */
            {8'h00}, /* 0x5db5 */
            {8'h00}, /* 0x5db4 */
            {8'h00}, /* 0x5db3 */
            {8'h00}, /* 0x5db2 */
            {8'h00}, /* 0x5db1 */
            {8'h00}, /* 0x5db0 */
            {8'h00}, /* 0x5daf */
            {8'h00}, /* 0x5dae */
            {8'h00}, /* 0x5dad */
            {8'h00}, /* 0x5dac */
            {8'h00}, /* 0x5dab */
            {8'h00}, /* 0x5daa */
            {8'h00}, /* 0x5da9 */
            {8'h00}, /* 0x5da8 */
            {8'h00}, /* 0x5da7 */
            {8'h00}, /* 0x5da6 */
            {8'h00}, /* 0x5da5 */
            {8'h00}, /* 0x5da4 */
            {8'h00}, /* 0x5da3 */
            {8'h00}, /* 0x5da2 */
            {8'h00}, /* 0x5da1 */
            {8'h00}, /* 0x5da0 */
            {8'h00}, /* 0x5d9f */
            {8'h00}, /* 0x5d9e */
            {8'h00}, /* 0x5d9d */
            {8'h00}, /* 0x5d9c */
            {8'h00}, /* 0x5d9b */
            {8'h00}, /* 0x5d9a */
            {8'h00}, /* 0x5d99 */
            {8'h00}, /* 0x5d98 */
            {8'h00}, /* 0x5d97 */
            {8'h00}, /* 0x5d96 */
            {8'h00}, /* 0x5d95 */
            {8'h00}, /* 0x5d94 */
            {8'h00}, /* 0x5d93 */
            {8'h00}, /* 0x5d92 */
            {8'h00}, /* 0x5d91 */
            {8'h00}, /* 0x5d90 */
            {8'h00}, /* 0x5d8f */
            {8'h00}, /* 0x5d8e */
            {8'h00}, /* 0x5d8d */
            {8'h00}, /* 0x5d8c */
            {8'h00}, /* 0x5d8b */
            {8'h00}, /* 0x5d8a */
            {8'h00}, /* 0x5d89 */
            {8'h00}, /* 0x5d88 */
            {8'h00}, /* 0x5d87 */
            {8'h00}, /* 0x5d86 */
            {8'h00}, /* 0x5d85 */
            {8'h00}, /* 0x5d84 */
            {8'h00}, /* 0x5d83 */
            {8'h00}, /* 0x5d82 */
            {8'h00}, /* 0x5d81 */
            {8'h00}, /* 0x5d80 */
            {8'h00}, /* 0x5d7f */
            {8'h00}, /* 0x5d7e */
            {8'h00}, /* 0x5d7d */
            {8'h00}, /* 0x5d7c */
            {8'h00}, /* 0x5d7b */
            {8'h00}, /* 0x5d7a */
            {8'h00}, /* 0x5d79 */
            {8'h00}, /* 0x5d78 */
            {8'h00}, /* 0x5d77 */
            {8'h00}, /* 0x5d76 */
            {8'h00}, /* 0x5d75 */
            {8'h00}, /* 0x5d74 */
            {8'h00}, /* 0x5d73 */
            {8'h00}, /* 0x5d72 */
            {8'h00}, /* 0x5d71 */
            {8'h00}, /* 0x5d70 */
            {8'h00}, /* 0x5d6f */
            {8'h00}, /* 0x5d6e */
            {8'h00}, /* 0x5d6d */
            {8'h00}, /* 0x5d6c */
            {8'h00}, /* 0x5d6b */
            {8'h00}, /* 0x5d6a */
            {8'h00}, /* 0x5d69 */
            {8'h00}, /* 0x5d68 */
            {8'h00}, /* 0x5d67 */
            {8'h00}, /* 0x5d66 */
            {8'h00}, /* 0x5d65 */
            {8'h00}, /* 0x5d64 */
            {8'h00}, /* 0x5d63 */
            {8'h00}, /* 0x5d62 */
            {8'h00}, /* 0x5d61 */
            {8'h00}, /* 0x5d60 */
            {8'h00}, /* 0x5d5f */
            {8'h00}, /* 0x5d5e */
            {8'h00}, /* 0x5d5d */
            {8'h00}, /* 0x5d5c */
            {8'h00}, /* 0x5d5b */
            {8'h00}, /* 0x5d5a */
            {8'h00}, /* 0x5d59 */
            {8'h00}, /* 0x5d58 */
            {8'h00}, /* 0x5d57 */
            {8'h00}, /* 0x5d56 */
            {8'h00}, /* 0x5d55 */
            {8'h00}, /* 0x5d54 */
            {8'h00}, /* 0x5d53 */
            {8'h00}, /* 0x5d52 */
            {8'h00}, /* 0x5d51 */
            {8'h00}, /* 0x5d50 */
            {8'h00}, /* 0x5d4f */
            {8'h00}, /* 0x5d4e */
            {8'h00}, /* 0x5d4d */
            {8'h00}, /* 0x5d4c */
            {8'h00}, /* 0x5d4b */
            {8'h00}, /* 0x5d4a */
            {8'h00}, /* 0x5d49 */
            {8'h00}, /* 0x5d48 */
            {8'h00}, /* 0x5d47 */
            {8'h00}, /* 0x5d46 */
            {8'h00}, /* 0x5d45 */
            {8'h00}, /* 0x5d44 */
            {8'h00}, /* 0x5d43 */
            {8'h00}, /* 0x5d42 */
            {8'h00}, /* 0x5d41 */
            {8'h00}, /* 0x5d40 */
            {8'h00}, /* 0x5d3f */
            {8'h00}, /* 0x5d3e */
            {8'h00}, /* 0x5d3d */
            {8'h00}, /* 0x5d3c */
            {8'h00}, /* 0x5d3b */
            {8'h00}, /* 0x5d3a */
            {8'h00}, /* 0x5d39 */
            {8'h00}, /* 0x5d38 */
            {8'h00}, /* 0x5d37 */
            {8'h00}, /* 0x5d36 */
            {8'h00}, /* 0x5d35 */
            {8'h00}, /* 0x5d34 */
            {8'h00}, /* 0x5d33 */
            {8'h00}, /* 0x5d32 */
            {8'h00}, /* 0x5d31 */
            {8'h00}, /* 0x5d30 */
            {8'h00}, /* 0x5d2f */
            {8'h00}, /* 0x5d2e */
            {8'h00}, /* 0x5d2d */
            {8'h00}, /* 0x5d2c */
            {8'h00}, /* 0x5d2b */
            {8'h00}, /* 0x5d2a */
            {8'h00}, /* 0x5d29 */
            {8'h00}, /* 0x5d28 */
            {8'h00}, /* 0x5d27 */
            {8'h00}, /* 0x5d26 */
            {8'h00}, /* 0x5d25 */
            {8'h00}, /* 0x5d24 */
            {8'h00}, /* 0x5d23 */
            {8'h00}, /* 0x5d22 */
            {8'h00}, /* 0x5d21 */
            {8'h00}, /* 0x5d20 */
            {8'h00}, /* 0x5d1f */
            {8'h00}, /* 0x5d1e */
            {8'h00}, /* 0x5d1d */
            {8'h00}, /* 0x5d1c */
            {8'h00}, /* 0x5d1b */
            {8'h00}, /* 0x5d1a */
            {8'h00}, /* 0x5d19 */
            {8'h00}, /* 0x5d18 */
            {8'h00}, /* 0x5d17 */
            {8'h00}, /* 0x5d16 */
            {8'h00}, /* 0x5d15 */
            {8'h00}, /* 0x5d14 */
            {8'h00}, /* 0x5d13 */
            {8'h00}, /* 0x5d12 */
            {8'h00}, /* 0x5d11 */
            {8'h00}, /* 0x5d10 */
            {8'h00}, /* 0x5d0f */
            {8'h00}, /* 0x5d0e */
            {8'h00}, /* 0x5d0d */
            {8'h00}, /* 0x5d0c */
            {8'h00}, /* 0x5d0b */
            {8'h00}, /* 0x5d0a */
            {8'h00}, /* 0x5d09 */
            {8'h00}, /* 0x5d08 */
            {8'h00}, /* 0x5d07 */
            {8'h00}, /* 0x5d06 */
            {8'h00}, /* 0x5d05 */
            {8'h00}, /* 0x5d04 */
            {8'h00}, /* 0x5d03 */
            {8'h00}, /* 0x5d02 */
            {8'h00}, /* 0x5d01 */
            {8'h00}, /* 0x5d00 */
            {8'h00}, /* 0x5cff */
            {8'h00}, /* 0x5cfe */
            {8'h00}, /* 0x5cfd */
            {8'h00}, /* 0x5cfc */
            {8'h00}, /* 0x5cfb */
            {8'h00}, /* 0x5cfa */
            {8'h00}, /* 0x5cf9 */
            {8'h00}, /* 0x5cf8 */
            {8'h00}, /* 0x5cf7 */
            {8'h00}, /* 0x5cf6 */
            {8'h00}, /* 0x5cf5 */
            {8'h00}, /* 0x5cf4 */
            {8'h00}, /* 0x5cf3 */
            {8'h00}, /* 0x5cf2 */
            {8'h00}, /* 0x5cf1 */
            {8'h00}, /* 0x5cf0 */
            {8'h00}, /* 0x5cef */
            {8'h00}, /* 0x5cee */
            {8'h00}, /* 0x5ced */
            {8'h00}, /* 0x5cec */
            {8'h00}, /* 0x5ceb */
            {8'h00}, /* 0x5cea */
            {8'h00}, /* 0x5ce9 */
            {8'h00}, /* 0x5ce8 */
            {8'h00}, /* 0x5ce7 */
            {8'h00}, /* 0x5ce6 */
            {8'h00}, /* 0x5ce5 */
            {8'h00}, /* 0x5ce4 */
            {8'h00}, /* 0x5ce3 */
            {8'h00}, /* 0x5ce2 */
            {8'h00}, /* 0x5ce1 */
            {8'h00}, /* 0x5ce0 */
            {8'h00}, /* 0x5cdf */
            {8'h00}, /* 0x5cde */
            {8'h00}, /* 0x5cdd */
            {8'h00}, /* 0x5cdc */
            {8'h00}, /* 0x5cdb */
            {8'h00}, /* 0x5cda */
            {8'h00}, /* 0x5cd9 */
            {8'h00}, /* 0x5cd8 */
            {8'h00}, /* 0x5cd7 */
            {8'h00}, /* 0x5cd6 */
            {8'h00}, /* 0x5cd5 */
            {8'h00}, /* 0x5cd4 */
            {8'h00}, /* 0x5cd3 */
            {8'h00}, /* 0x5cd2 */
            {8'h00}, /* 0x5cd1 */
            {8'h00}, /* 0x5cd0 */
            {8'h00}, /* 0x5ccf */
            {8'h00}, /* 0x5cce */
            {8'h00}, /* 0x5ccd */
            {8'h00}, /* 0x5ccc */
            {8'h00}, /* 0x5ccb */
            {8'h00}, /* 0x5cca */
            {8'h00}, /* 0x5cc9 */
            {8'h00}, /* 0x5cc8 */
            {8'h00}, /* 0x5cc7 */
            {8'h00}, /* 0x5cc6 */
            {8'h00}, /* 0x5cc5 */
            {8'h00}, /* 0x5cc4 */
            {8'h00}, /* 0x5cc3 */
            {8'h00}, /* 0x5cc2 */
            {8'h00}, /* 0x5cc1 */
            {8'h00}, /* 0x5cc0 */
            {8'h00}, /* 0x5cbf */
            {8'h00}, /* 0x5cbe */
            {8'h00}, /* 0x5cbd */
            {8'h00}, /* 0x5cbc */
            {8'h00}, /* 0x5cbb */
            {8'h00}, /* 0x5cba */
            {8'h00}, /* 0x5cb9 */
            {8'h00}, /* 0x5cb8 */
            {8'h00}, /* 0x5cb7 */
            {8'h00}, /* 0x5cb6 */
            {8'h00}, /* 0x5cb5 */
            {8'h00}, /* 0x5cb4 */
            {8'h00}, /* 0x5cb3 */
            {8'h00}, /* 0x5cb2 */
            {8'h00}, /* 0x5cb1 */
            {8'h00}, /* 0x5cb0 */
            {8'h00}, /* 0x5caf */
            {8'h00}, /* 0x5cae */
            {8'h00}, /* 0x5cad */
            {8'h00}, /* 0x5cac */
            {8'h00}, /* 0x5cab */
            {8'h00}, /* 0x5caa */
            {8'h00}, /* 0x5ca9 */
            {8'h00}, /* 0x5ca8 */
            {8'h00}, /* 0x5ca7 */
            {8'h00}, /* 0x5ca6 */
            {8'h00}, /* 0x5ca5 */
            {8'h00}, /* 0x5ca4 */
            {8'h00}, /* 0x5ca3 */
            {8'h00}, /* 0x5ca2 */
            {8'h00}, /* 0x5ca1 */
            {8'h00}, /* 0x5ca0 */
            {8'h00}, /* 0x5c9f */
            {8'h00}, /* 0x5c9e */
            {8'h00}, /* 0x5c9d */
            {8'h00}, /* 0x5c9c */
            {8'h00}, /* 0x5c9b */
            {8'h00}, /* 0x5c9a */
            {8'h00}, /* 0x5c99 */
            {8'h00}, /* 0x5c98 */
            {8'h00}, /* 0x5c97 */
            {8'h00}, /* 0x5c96 */
            {8'h00}, /* 0x5c95 */
            {8'h00}, /* 0x5c94 */
            {8'h00}, /* 0x5c93 */
            {8'h00}, /* 0x5c92 */
            {8'h00}, /* 0x5c91 */
            {8'h00}, /* 0x5c90 */
            {8'h00}, /* 0x5c8f */
            {8'h00}, /* 0x5c8e */
            {8'h00}, /* 0x5c8d */
            {8'h00}, /* 0x5c8c */
            {8'h00}, /* 0x5c8b */
            {8'h00}, /* 0x5c8a */
            {8'h00}, /* 0x5c89 */
            {8'h00}, /* 0x5c88 */
            {8'h00}, /* 0x5c87 */
            {8'h00}, /* 0x5c86 */
            {8'h00}, /* 0x5c85 */
            {8'h00}, /* 0x5c84 */
            {8'h00}, /* 0x5c83 */
            {8'h00}, /* 0x5c82 */
            {8'h00}, /* 0x5c81 */
            {8'h00}, /* 0x5c80 */
            {8'h00}, /* 0x5c7f */
            {8'h00}, /* 0x5c7e */
            {8'h00}, /* 0x5c7d */
            {8'h00}, /* 0x5c7c */
            {8'h00}, /* 0x5c7b */
            {8'h00}, /* 0x5c7a */
            {8'h00}, /* 0x5c79 */
            {8'h00}, /* 0x5c78 */
            {8'h00}, /* 0x5c77 */
            {8'h00}, /* 0x5c76 */
            {8'h00}, /* 0x5c75 */
            {8'h00}, /* 0x5c74 */
            {8'h00}, /* 0x5c73 */
            {8'h00}, /* 0x5c72 */
            {8'h00}, /* 0x5c71 */
            {8'h00}, /* 0x5c70 */
            {8'h00}, /* 0x5c6f */
            {8'h00}, /* 0x5c6e */
            {8'h00}, /* 0x5c6d */
            {8'h00}, /* 0x5c6c */
            {8'h00}, /* 0x5c6b */
            {8'h00}, /* 0x5c6a */
            {8'h00}, /* 0x5c69 */
            {8'h00}, /* 0x5c68 */
            {8'h00}, /* 0x5c67 */
            {8'h00}, /* 0x5c66 */
            {8'h00}, /* 0x5c65 */
            {8'h00}, /* 0x5c64 */
            {8'h00}, /* 0x5c63 */
            {8'h00}, /* 0x5c62 */
            {8'h00}, /* 0x5c61 */
            {8'h00}, /* 0x5c60 */
            {8'h00}, /* 0x5c5f */
            {8'h00}, /* 0x5c5e */
            {8'h00}, /* 0x5c5d */
            {8'h00}, /* 0x5c5c */
            {8'h00}, /* 0x5c5b */
            {8'h00}, /* 0x5c5a */
            {8'h00}, /* 0x5c59 */
            {8'h00}, /* 0x5c58 */
            {8'h00}, /* 0x5c57 */
            {8'h00}, /* 0x5c56 */
            {8'h00}, /* 0x5c55 */
            {8'h00}, /* 0x5c54 */
            {8'h00}, /* 0x5c53 */
            {8'h00}, /* 0x5c52 */
            {8'h00}, /* 0x5c51 */
            {8'h00}, /* 0x5c50 */
            {8'h00}, /* 0x5c4f */
            {8'h00}, /* 0x5c4e */
            {8'h00}, /* 0x5c4d */
            {8'h00}, /* 0x5c4c */
            {8'h00}, /* 0x5c4b */
            {8'h00}, /* 0x5c4a */
            {8'h00}, /* 0x5c49 */
            {8'h00}, /* 0x5c48 */
            {8'h00}, /* 0x5c47 */
            {8'h00}, /* 0x5c46 */
            {8'h00}, /* 0x5c45 */
            {8'h00}, /* 0x5c44 */
            {8'h00}, /* 0x5c43 */
            {8'h00}, /* 0x5c42 */
            {8'h00}, /* 0x5c41 */
            {8'h00}, /* 0x5c40 */
            {8'h00}, /* 0x5c3f */
            {8'h00}, /* 0x5c3e */
            {8'h00}, /* 0x5c3d */
            {8'h00}, /* 0x5c3c */
            {8'h00}, /* 0x5c3b */
            {8'h00}, /* 0x5c3a */
            {8'h00}, /* 0x5c39 */
            {8'h00}, /* 0x5c38 */
            {8'h00}, /* 0x5c37 */
            {8'h00}, /* 0x5c36 */
            {8'h00}, /* 0x5c35 */
            {8'h00}, /* 0x5c34 */
            {8'h00}, /* 0x5c33 */
            {8'h00}, /* 0x5c32 */
            {8'h00}, /* 0x5c31 */
            {8'h00}, /* 0x5c30 */
            {8'h00}, /* 0x5c2f */
            {8'h00}, /* 0x5c2e */
            {8'h00}, /* 0x5c2d */
            {8'h00}, /* 0x5c2c */
            {8'h00}, /* 0x5c2b */
            {8'h00}, /* 0x5c2a */
            {8'h00}, /* 0x5c29 */
            {8'h00}, /* 0x5c28 */
            {8'h00}, /* 0x5c27 */
            {8'h00}, /* 0x5c26 */
            {8'h00}, /* 0x5c25 */
            {8'h00}, /* 0x5c24 */
            {8'h00}, /* 0x5c23 */
            {8'h00}, /* 0x5c22 */
            {8'h00}, /* 0x5c21 */
            {8'h00}, /* 0x5c20 */
            {8'h00}, /* 0x5c1f */
            {8'h00}, /* 0x5c1e */
            {8'h00}, /* 0x5c1d */
            {8'h00}, /* 0x5c1c */
            {8'h00}, /* 0x5c1b */
            {8'h00}, /* 0x5c1a */
            {8'h00}, /* 0x5c19 */
            {8'h00}, /* 0x5c18 */
            {8'h00}, /* 0x5c17 */
            {8'h00}, /* 0x5c16 */
            {8'h00}, /* 0x5c15 */
            {8'h00}, /* 0x5c14 */
            {8'h00}, /* 0x5c13 */
            {8'h00}, /* 0x5c12 */
            {8'h00}, /* 0x5c11 */
            {8'h00}, /* 0x5c10 */
            {8'h00}, /* 0x5c0f */
            {8'h00}, /* 0x5c0e */
            {8'h00}, /* 0x5c0d */
            {8'h00}, /* 0x5c0c */
            {8'h00}, /* 0x5c0b */
            {8'h00}, /* 0x5c0a */
            {8'h00}, /* 0x5c09 */
            {8'h00}, /* 0x5c08 */
            {8'h00}, /* 0x5c07 */
            {8'h00}, /* 0x5c06 */
            {8'h00}, /* 0x5c05 */
            {8'h00}, /* 0x5c04 */
            {8'h00}, /* 0x5c03 */
            {8'h00}, /* 0x5c02 */
            {8'h00}, /* 0x5c01 */
            {8'h00}, /* 0x5c00 */
            {8'h00}, /* 0x5bff */
            {8'h00}, /* 0x5bfe */
            {8'h00}, /* 0x5bfd */
            {8'h00}, /* 0x5bfc */
            {8'h00}, /* 0x5bfb */
            {8'h00}, /* 0x5bfa */
            {8'h00}, /* 0x5bf9 */
            {8'h00}, /* 0x5bf8 */
            {8'h00}, /* 0x5bf7 */
            {8'h00}, /* 0x5bf6 */
            {8'h00}, /* 0x5bf5 */
            {8'h00}, /* 0x5bf4 */
            {8'h00}, /* 0x5bf3 */
            {8'h00}, /* 0x5bf2 */
            {8'h00}, /* 0x5bf1 */
            {8'h00}, /* 0x5bf0 */
            {8'h00}, /* 0x5bef */
            {8'h00}, /* 0x5bee */
            {8'h00}, /* 0x5bed */
            {8'h00}, /* 0x5bec */
            {8'h00}, /* 0x5beb */
            {8'h00}, /* 0x5bea */
            {8'h00}, /* 0x5be9 */
            {8'h00}, /* 0x5be8 */
            {8'h00}, /* 0x5be7 */
            {8'h00}, /* 0x5be6 */
            {8'h00}, /* 0x5be5 */
            {8'h00}, /* 0x5be4 */
            {8'h00}, /* 0x5be3 */
            {8'h00}, /* 0x5be2 */
            {8'h00}, /* 0x5be1 */
            {8'h00}, /* 0x5be0 */
            {8'h00}, /* 0x5bdf */
            {8'h00}, /* 0x5bde */
            {8'h00}, /* 0x5bdd */
            {8'h00}, /* 0x5bdc */
            {8'h00}, /* 0x5bdb */
            {8'h00}, /* 0x5bda */
            {8'h00}, /* 0x5bd9 */
            {8'h00}, /* 0x5bd8 */
            {8'h00}, /* 0x5bd7 */
            {8'h00}, /* 0x5bd6 */
            {8'h00}, /* 0x5bd5 */
            {8'h00}, /* 0x5bd4 */
            {8'h00}, /* 0x5bd3 */
            {8'h00}, /* 0x5bd2 */
            {8'h00}, /* 0x5bd1 */
            {8'h00}, /* 0x5bd0 */
            {8'h00}, /* 0x5bcf */
            {8'h00}, /* 0x5bce */
            {8'h00}, /* 0x5bcd */
            {8'h00}, /* 0x5bcc */
            {8'h00}, /* 0x5bcb */
            {8'h00}, /* 0x5bca */
            {8'h00}, /* 0x5bc9 */
            {8'h00}, /* 0x5bc8 */
            {8'h00}, /* 0x5bc7 */
            {8'h00}, /* 0x5bc6 */
            {8'h00}, /* 0x5bc5 */
            {8'h00}, /* 0x5bc4 */
            {8'h00}, /* 0x5bc3 */
            {8'h00}, /* 0x5bc2 */
            {8'h00}, /* 0x5bc1 */
            {8'h00}, /* 0x5bc0 */
            {8'h00}, /* 0x5bbf */
            {8'h00}, /* 0x5bbe */
            {8'h00}, /* 0x5bbd */
            {8'h00}, /* 0x5bbc */
            {8'h00}, /* 0x5bbb */
            {8'h00}, /* 0x5bba */
            {8'h00}, /* 0x5bb9 */
            {8'h00}, /* 0x5bb8 */
            {8'h00}, /* 0x5bb7 */
            {8'h00}, /* 0x5bb6 */
            {8'h00}, /* 0x5bb5 */
            {8'h00}, /* 0x5bb4 */
            {8'h00}, /* 0x5bb3 */
            {8'h00}, /* 0x5bb2 */
            {8'h00}, /* 0x5bb1 */
            {8'h00}, /* 0x5bb0 */
            {8'h00}, /* 0x5baf */
            {8'h00}, /* 0x5bae */
            {8'h00}, /* 0x5bad */
            {8'h00}, /* 0x5bac */
            {8'h00}, /* 0x5bab */
            {8'h00}, /* 0x5baa */
            {8'h00}, /* 0x5ba9 */
            {8'h00}, /* 0x5ba8 */
            {8'h00}, /* 0x5ba7 */
            {8'h00}, /* 0x5ba6 */
            {8'h00}, /* 0x5ba5 */
            {8'h00}, /* 0x5ba4 */
            {8'h00}, /* 0x5ba3 */
            {8'h00}, /* 0x5ba2 */
            {8'h00}, /* 0x5ba1 */
            {8'h00}, /* 0x5ba0 */
            {8'h00}, /* 0x5b9f */
            {8'h00}, /* 0x5b9e */
            {8'h00}, /* 0x5b9d */
            {8'h00}, /* 0x5b9c */
            {8'h00}, /* 0x5b9b */
            {8'h00}, /* 0x5b9a */
            {8'h00}, /* 0x5b99 */
            {8'h00}, /* 0x5b98 */
            {8'h00}, /* 0x5b97 */
            {8'h00}, /* 0x5b96 */
            {8'h00}, /* 0x5b95 */
            {8'h00}, /* 0x5b94 */
            {8'h00}, /* 0x5b93 */
            {8'h00}, /* 0x5b92 */
            {8'h00}, /* 0x5b91 */
            {8'h00}, /* 0x5b90 */
            {8'h00}, /* 0x5b8f */
            {8'h00}, /* 0x5b8e */
            {8'h00}, /* 0x5b8d */
            {8'h00}, /* 0x5b8c */
            {8'h00}, /* 0x5b8b */
            {8'h00}, /* 0x5b8a */
            {8'h00}, /* 0x5b89 */
            {8'h00}, /* 0x5b88 */
            {8'h00}, /* 0x5b87 */
            {8'h00}, /* 0x5b86 */
            {8'h00}, /* 0x5b85 */
            {8'h00}, /* 0x5b84 */
            {8'h00}, /* 0x5b83 */
            {8'h00}, /* 0x5b82 */
            {8'h00}, /* 0x5b81 */
            {8'h00}, /* 0x5b80 */
            {8'h00}, /* 0x5b7f */
            {8'h00}, /* 0x5b7e */
            {8'h00}, /* 0x5b7d */
            {8'h00}, /* 0x5b7c */
            {8'h00}, /* 0x5b7b */
            {8'h00}, /* 0x5b7a */
            {8'h00}, /* 0x5b79 */
            {8'h00}, /* 0x5b78 */
            {8'h00}, /* 0x5b77 */
            {8'h00}, /* 0x5b76 */
            {8'h00}, /* 0x5b75 */
            {8'h00}, /* 0x5b74 */
            {8'h00}, /* 0x5b73 */
            {8'h00}, /* 0x5b72 */
            {8'h00}, /* 0x5b71 */
            {8'h00}, /* 0x5b70 */
            {8'h00}, /* 0x5b6f */
            {8'h00}, /* 0x5b6e */
            {8'h00}, /* 0x5b6d */
            {8'h00}, /* 0x5b6c */
            {8'h00}, /* 0x5b6b */
            {8'h00}, /* 0x5b6a */
            {8'h00}, /* 0x5b69 */
            {8'h00}, /* 0x5b68 */
            {8'h00}, /* 0x5b67 */
            {8'h00}, /* 0x5b66 */
            {8'h00}, /* 0x5b65 */
            {8'h00}, /* 0x5b64 */
            {8'h00}, /* 0x5b63 */
            {8'h00}, /* 0x5b62 */
            {8'h00}, /* 0x5b61 */
            {8'h00}, /* 0x5b60 */
            {8'h00}, /* 0x5b5f */
            {8'h00}, /* 0x5b5e */
            {8'h00}, /* 0x5b5d */
            {8'h00}, /* 0x5b5c */
            {8'h00}, /* 0x5b5b */
            {8'h00}, /* 0x5b5a */
            {8'h00}, /* 0x5b59 */
            {8'h00}, /* 0x5b58 */
            {8'h00}, /* 0x5b57 */
            {8'h00}, /* 0x5b56 */
            {8'h00}, /* 0x5b55 */
            {8'h00}, /* 0x5b54 */
            {8'h00}, /* 0x5b53 */
            {8'h00}, /* 0x5b52 */
            {8'h00}, /* 0x5b51 */
            {8'h00}, /* 0x5b50 */
            {8'h00}, /* 0x5b4f */
            {8'h00}, /* 0x5b4e */
            {8'h00}, /* 0x5b4d */
            {8'h00}, /* 0x5b4c */
            {8'h00}, /* 0x5b4b */
            {8'h00}, /* 0x5b4a */
            {8'h00}, /* 0x5b49 */
            {8'h00}, /* 0x5b48 */
            {8'h00}, /* 0x5b47 */
            {8'h00}, /* 0x5b46 */
            {8'h00}, /* 0x5b45 */
            {8'h00}, /* 0x5b44 */
            {8'h00}, /* 0x5b43 */
            {8'h00}, /* 0x5b42 */
            {8'h00}, /* 0x5b41 */
            {8'h00}, /* 0x5b40 */
            {8'h00}, /* 0x5b3f */
            {8'h00}, /* 0x5b3e */
            {8'h00}, /* 0x5b3d */
            {8'h00}, /* 0x5b3c */
            {8'h00}, /* 0x5b3b */
            {8'h00}, /* 0x5b3a */
            {8'h00}, /* 0x5b39 */
            {8'h00}, /* 0x5b38 */
            {8'h00}, /* 0x5b37 */
            {8'h00}, /* 0x5b36 */
            {8'h00}, /* 0x5b35 */
            {8'h00}, /* 0x5b34 */
            {8'h00}, /* 0x5b33 */
            {8'h00}, /* 0x5b32 */
            {8'h00}, /* 0x5b31 */
            {8'h00}, /* 0x5b30 */
            {8'h00}, /* 0x5b2f */
            {8'h00}, /* 0x5b2e */
            {8'h00}, /* 0x5b2d */
            {8'h00}, /* 0x5b2c */
            {8'h00}, /* 0x5b2b */
            {8'h00}, /* 0x5b2a */
            {8'h00}, /* 0x5b29 */
            {8'h00}, /* 0x5b28 */
            {8'h00}, /* 0x5b27 */
            {8'h00}, /* 0x5b26 */
            {8'h00}, /* 0x5b25 */
            {8'h00}, /* 0x5b24 */
            {8'h00}, /* 0x5b23 */
            {8'h00}, /* 0x5b22 */
            {8'h00}, /* 0x5b21 */
            {8'h00}, /* 0x5b20 */
            {8'h00}, /* 0x5b1f */
            {8'h00}, /* 0x5b1e */
            {8'h00}, /* 0x5b1d */
            {8'h00}, /* 0x5b1c */
            {8'h00}, /* 0x5b1b */
            {8'h00}, /* 0x5b1a */
            {8'h00}, /* 0x5b19 */
            {8'h00}, /* 0x5b18 */
            {8'h00}, /* 0x5b17 */
            {8'h00}, /* 0x5b16 */
            {8'h00}, /* 0x5b15 */
            {8'h00}, /* 0x5b14 */
            {8'h00}, /* 0x5b13 */
            {8'h00}, /* 0x5b12 */
            {8'h00}, /* 0x5b11 */
            {8'h00}, /* 0x5b10 */
            {8'h00}, /* 0x5b0f */
            {8'h00}, /* 0x5b0e */
            {8'h00}, /* 0x5b0d */
            {8'h00}, /* 0x5b0c */
            {8'h00}, /* 0x5b0b */
            {8'h00}, /* 0x5b0a */
            {8'h00}, /* 0x5b09 */
            {8'h00}, /* 0x5b08 */
            {8'h00}, /* 0x5b07 */
            {8'h00}, /* 0x5b06 */
            {8'h00}, /* 0x5b05 */
            {8'h00}, /* 0x5b04 */
            {8'h00}, /* 0x5b03 */
            {8'h00}, /* 0x5b02 */
            {8'h00}, /* 0x5b01 */
            {8'h00}, /* 0x5b00 */
            {8'h00}, /* 0x5aff */
            {8'h00}, /* 0x5afe */
            {8'h00}, /* 0x5afd */
            {8'h00}, /* 0x5afc */
            {8'h00}, /* 0x5afb */
            {8'h00}, /* 0x5afa */
            {8'h00}, /* 0x5af9 */
            {8'h00}, /* 0x5af8 */
            {8'h00}, /* 0x5af7 */
            {8'h00}, /* 0x5af6 */
            {8'h00}, /* 0x5af5 */
            {8'h00}, /* 0x5af4 */
            {8'h00}, /* 0x5af3 */
            {8'h00}, /* 0x5af2 */
            {8'h00}, /* 0x5af1 */
            {8'h00}, /* 0x5af0 */
            {8'h00}, /* 0x5aef */
            {8'h00}, /* 0x5aee */
            {8'h00}, /* 0x5aed */
            {8'h00}, /* 0x5aec */
            {8'h00}, /* 0x5aeb */
            {8'h00}, /* 0x5aea */
            {8'h00}, /* 0x5ae9 */
            {8'h00}, /* 0x5ae8 */
            {8'h00}, /* 0x5ae7 */
            {8'h00}, /* 0x5ae6 */
            {8'h00}, /* 0x5ae5 */
            {8'h00}, /* 0x5ae4 */
            {8'h00}, /* 0x5ae3 */
            {8'h00}, /* 0x5ae2 */
            {8'h00}, /* 0x5ae1 */
            {8'h00}, /* 0x5ae0 */
            {8'h00}, /* 0x5adf */
            {8'h00}, /* 0x5ade */
            {8'h00}, /* 0x5add */
            {8'h00}, /* 0x5adc */
            {8'h00}, /* 0x5adb */
            {8'h00}, /* 0x5ada */
            {8'h00}, /* 0x5ad9 */
            {8'h00}, /* 0x5ad8 */
            {8'h00}, /* 0x5ad7 */
            {8'h00}, /* 0x5ad6 */
            {8'h00}, /* 0x5ad5 */
            {8'h00}, /* 0x5ad4 */
            {8'h00}, /* 0x5ad3 */
            {8'h00}, /* 0x5ad2 */
            {8'h00}, /* 0x5ad1 */
            {8'h00}, /* 0x5ad0 */
            {8'h00}, /* 0x5acf */
            {8'h00}, /* 0x5ace */
            {8'h00}, /* 0x5acd */
            {8'h00}, /* 0x5acc */
            {8'h00}, /* 0x5acb */
            {8'h00}, /* 0x5aca */
            {8'h00}, /* 0x5ac9 */
            {8'h00}, /* 0x5ac8 */
            {8'h00}, /* 0x5ac7 */
            {8'h00}, /* 0x5ac6 */
            {8'h00}, /* 0x5ac5 */
            {8'h00}, /* 0x5ac4 */
            {8'h00}, /* 0x5ac3 */
            {8'h00}, /* 0x5ac2 */
            {8'h00}, /* 0x5ac1 */
            {8'h00}, /* 0x5ac0 */
            {8'h00}, /* 0x5abf */
            {8'h00}, /* 0x5abe */
            {8'h00}, /* 0x5abd */
            {8'h00}, /* 0x5abc */
            {8'h00}, /* 0x5abb */
            {8'h00}, /* 0x5aba */
            {8'h00}, /* 0x5ab9 */
            {8'h00}, /* 0x5ab8 */
            {8'h00}, /* 0x5ab7 */
            {8'h00}, /* 0x5ab6 */
            {8'h00}, /* 0x5ab5 */
            {8'h00}, /* 0x5ab4 */
            {8'h00}, /* 0x5ab3 */
            {8'h00}, /* 0x5ab2 */
            {8'h00}, /* 0x5ab1 */
            {8'h00}, /* 0x5ab0 */
            {8'h00}, /* 0x5aaf */
            {8'h00}, /* 0x5aae */
            {8'h00}, /* 0x5aad */
            {8'h00}, /* 0x5aac */
            {8'h00}, /* 0x5aab */
            {8'h00}, /* 0x5aaa */
            {8'h00}, /* 0x5aa9 */
            {8'h00}, /* 0x5aa8 */
            {8'h00}, /* 0x5aa7 */
            {8'h00}, /* 0x5aa6 */
            {8'h00}, /* 0x5aa5 */
            {8'h00}, /* 0x5aa4 */
            {8'h00}, /* 0x5aa3 */
            {8'h00}, /* 0x5aa2 */
            {8'h00}, /* 0x5aa1 */
            {8'h00}, /* 0x5aa0 */
            {8'h00}, /* 0x5a9f */
            {8'h00}, /* 0x5a9e */
            {8'h00}, /* 0x5a9d */
            {8'h00}, /* 0x5a9c */
            {8'h00}, /* 0x5a9b */
            {8'h00}, /* 0x5a9a */
            {8'h00}, /* 0x5a99 */
            {8'h00}, /* 0x5a98 */
            {8'h00}, /* 0x5a97 */
            {8'h00}, /* 0x5a96 */
            {8'h00}, /* 0x5a95 */
            {8'h00}, /* 0x5a94 */
            {8'h00}, /* 0x5a93 */
            {8'h00}, /* 0x5a92 */
            {8'h00}, /* 0x5a91 */
            {8'h00}, /* 0x5a90 */
            {8'h00}, /* 0x5a8f */
            {8'h00}, /* 0x5a8e */
            {8'h00}, /* 0x5a8d */
            {8'h00}, /* 0x5a8c */
            {8'h00}, /* 0x5a8b */
            {8'h00}, /* 0x5a8a */
            {8'h00}, /* 0x5a89 */
            {8'h00}, /* 0x5a88 */
            {8'h00}, /* 0x5a87 */
            {8'h00}, /* 0x5a86 */
            {8'h00}, /* 0x5a85 */
            {8'h00}, /* 0x5a84 */
            {8'h00}, /* 0x5a83 */
            {8'h00}, /* 0x5a82 */
            {8'h00}, /* 0x5a81 */
            {8'h00}, /* 0x5a80 */
            {8'h00}, /* 0x5a7f */
            {8'h00}, /* 0x5a7e */
            {8'h00}, /* 0x5a7d */
            {8'h00}, /* 0x5a7c */
            {8'h00}, /* 0x5a7b */
            {8'h00}, /* 0x5a7a */
            {8'h00}, /* 0x5a79 */
            {8'h00}, /* 0x5a78 */
            {8'h00}, /* 0x5a77 */
            {8'h00}, /* 0x5a76 */
            {8'h00}, /* 0x5a75 */
            {8'h00}, /* 0x5a74 */
            {8'h00}, /* 0x5a73 */
            {8'h00}, /* 0x5a72 */
            {8'h00}, /* 0x5a71 */
            {8'h00}, /* 0x5a70 */
            {8'h00}, /* 0x5a6f */
            {8'h00}, /* 0x5a6e */
            {8'h00}, /* 0x5a6d */
            {8'h00}, /* 0x5a6c */
            {8'h00}, /* 0x5a6b */
            {8'h00}, /* 0x5a6a */
            {8'h00}, /* 0x5a69 */
            {8'h00}, /* 0x5a68 */
            {8'h00}, /* 0x5a67 */
            {8'h00}, /* 0x5a66 */
            {8'h00}, /* 0x5a65 */
            {8'h00}, /* 0x5a64 */
            {8'h00}, /* 0x5a63 */
            {8'h00}, /* 0x5a62 */
            {8'h00}, /* 0x5a61 */
            {8'h00}, /* 0x5a60 */
            {8'h00}, /* 0x5a5f */
            {8'h00}, /* 0x5a5e */
            {8'h00}, /* 0x5a5d */
            {8'h00}, /* 0x5a5c */
            {8'h00}, /* 0x5a5b */
            {8'h00}, /* 0x5a5a */
            {8'h00}, /* 0x5a59 */
            {8'h00}, /* 0x5a58 */
            {8'h00}, /* 0x5a57 */
            {8'h00}, /* 0x5a56 */
            {8'h00}, /* 0x5a55 */
            {8'h00}, /* 0x5a54 */
            {8'h00}, /* 0x5a53 */
            {8'h00}, /* 0x5a52 */
            {8'h00}, /* 0x5a51 */
            {8'h00}, /* 0x5a50 */
            {8'h00}, /* 0x5a4f */
            {8'h00}, /* 0x5a4e */
            {8'h00}, /* 0x5a4d */
            {8'h00}, /* 0x5a4c */
            {8'h00}, /* 0x5a4b */
            {8'h00}, /* 0x5a4a */
            {8'h00}, /* 0x5a49 */
            {8'h00}, /* 0x5a48 */
            {8'h00}, /* 0x5a47 */
            {8'h00}, /* 0x5a46 */
            {8'h00}, /* 0x5a45 */
            {8'h00}, /* 0x5a44 */
            {8'h00}, /* 0x5a43 */
            {8'h00}, /* 0x5a42 */
            {8'h00}, /* 0x5a41 */
            {8'h00}, /* 0x5a40 */
            {8'h00}, /* 0x5a3f */
            {8'h00}, /* 0x5a3e */
            {8'h00}, /* 0x5a3d */
            {8'h00}, /* 0x5a3c */
            {8'h00}, /* 0x5a3b */
            {8'h00}, /* 0x5a3a */
            {8'h00}, /* 0x5a39 */
            {8'h00}, /* 0x5a38 */
            {8'h00}, /* 0x5a37 */
            {8'h00}, /* 0x5a36 */
            {8'h00}, /* 0x5a35 */
            {8'h00}, /* 0x5a34 */
            {8'h00}, /* 0x5a33 */
            {8'h00}, /* 0x5a32 */
            {8'h00}, /* 0x5a31 */
            {8'h00}, /* 0x5a30 */
            {8'h00}, /* 0x5a2f */
            {8'h00}, /* 0x5a2e */
            {8'h00}, /* 0x5a2d */
            {8'h00}, /* 0x5a2c */
            {8'h00}, /* 0x5a2b */
            {8'h00}, /* 0x5a2a */
            {8'h00}, /* 0x5a29 */
            {8'h00}, /* 0x5a28 */
            {8'h00}, /* 0x5a27 */
            {8'h00}, /* 0x5a26 */
            {8'h00}, /* 0x5a25 */
            {8'h00}, /* 0x5a24 */
            {8'h00}, /* 0x5a23 */
            {8'h00}, /* 0x5a22 */
            {8'h00}, /* 0x5a21 */
            {8'h00}, /* 0x5a20 */
            {8'h00}, /* 0x5a1f */
            {8'h00}, /* 0x5a1e */
            {8'h00}, /* 0x5a1d */
            {8'h00}, /* 0x5a1c */
            {8'h00}, /* 0x5a1b */
            {8'h00}, /* 0x5a1a */
            {8'h00}, /* 0x5a19 */
            {8'h00}, /* 0x5a18 */
            {8'h00}, /* 0x5a17 */
            {8'h00}, /* 0x5a16 */
            {8'h00}, /* 0x5a15 */
            {8'h00}, /* 0x5a14 */
            {8'h00}, /* 0x5a13 */
            {8'h00}, /* 0x5a12 */
            {8'h00}, /* 0x5a11 */
            {8'h00}, /* 0x5a10 */
            {8'h00}, /* 0x5a0f */
            {8'h00}, /* 0x5a0e */
            {8'h00}, /* 0x5a0d */
            {8'h00}, /* 0x5a0c */
            {8'h00}, /* 0x5a0b */
            {8'h00}, /* 0x5a0a */
            {8'h00}, /* 0x5a09 */
            {8'h00}, /* 0x5a08 */
            {8'h00}, /* 0x5a07 */
            {8'h00}, /* 0x5a06 */
            {8'h00}, /* 0x5a05 */
            {8'h00}, /* 0x5a04 */
            {8'h00}, /* 0x5a03 */
            {8'h00}, /* 0x5a02 */
            {8'h00}, /* 0x5a01 */
            {8'h00}, /* 0x5a00 */
            {8'h00}, /* 0x59ff */
            {8'h00}, /* 0x59fe */
            {8'h00}, /* 0x59fd */
            {8'h00}, /* 0x59fc */
            {8'h00}, /* 0x59fb */
            {8'h00}, /* 0x59fa */
            {8'h00}, /* 0x59f9 */
            {8'h00}, /* 0x59f8 */
            {8'h00}, /* 0x59f7 */
            {8'h00}, /* 0x59f6 */
            {8'h00}, /* 0x59f5 */
            {8'h00}, /* 0x59f4 */
            {8'h00}, /* 0x59f3 */
            {8'h00}, /* 0x59f2 */
            {8'h00}, /* 0x59f1 */
            {8'h00}, /* 0x59f0 */
            {8'h00}, /* 0x59ef */
            {8'h00}, /* 0x59ee */
            {8'h00}, /* 0x59ed */
            {8'h00}, /* 0x59ec */
            {8'h00}, /* 0x59eb */
            {8'h00}, /* 0x59ea */
            {8'h00}, /* 0x59e9 */
            {8'h00}, /* 0x59e8 */
            {8'h00}, /* 0x59e7 */
            {8'h00}, /* 0x59e6 */
            {8'h00}, /* 0x59e5 */
            {8'h00}, /* 0x59e4 */
            {8'h00}, /* 0x59e3 */
            {8'h00}, /* 0x59e2 */
            {8'h00}, /* 0x59e1 */
            {8'h00}, /* 0x59e0 */
            {8'h00}, /* 0x59df */
            {8'h00}, /* 0x59de */
            {8'h00}, /* 0x59dd */
            {8'h00}, /* 0x59dc */
            {8'h00}, /* 0x59db */
            {8'h00}, /* 0x59da */
            {8'h00}, /* 0x59d9 */
            {8'h00}, /* 0x59d8 */
            {8'h00}, /* 0x59d7 */
            {8'h00}, /* 0x59d6 */
            {8'h00}, /* 0x59d5 */
            {8'h00}, /* 0x59d4 */
            {8'h00}, /* 0x59d3 */
            {8'h00}, /* 0x59d2 */
            {8'h00}, /* 0x59d1 */
            {8'h00}, /* 0x59d0 */
            {8'h00}, /* 0x59cf */
            {8'h00}, /* 0x59ce */
            {8'h00}, /* 0x59cd */
            {8'h00}, /* 0x59cc */
            {8'h00}, /* 0x59cb */
            {8'h00}, /* 0x59ca */
            {8'h00}, /* 0x59c9 */
            {8'h00}, /* 0x59c8 */
            {8'h00}, /* 0x59c7 */
            {8'h00}, /* 0x59c6 */
            {8'h00}, /* 0x59c5 */
            {8'h00}, /* 0x59c4 */
            {8'h00}, /* 0x59c3 */
            {8'h00}, /* 0x59c2 */
            {8'h00}, /* 0x59c1 */
            {8'h00}, /* 0x59c0 */
            {8'h00}, /* 0x59bf */
            {8'h00}, /* 0x59be */
            {8'h00}, /* 0x59bd */
            {8'h00}, /* 0x59bc */
            {8'h00}, /* 0x59bb */
            {8'h00}, /* 0x59ba */
            {8'h00}, /* 0x59b9 */
            {8'h00}, /* 0x59b8 */
            {8'h00}, /* 0x59b7 */
            {8'h00}, /* 0x59b6 */
            {8'h00}, /* 0x59b5 */
            {8'h00}, /* 0x59b4 */
            {8'h00}, /* 0x59b3 */
            {8'h00}, /* 0x59b2 */
            {8'h00}, /* 0x59b1 */
            {8'h00}, /* 0x59b0 */
            {8'h00}, /* 0x59af */
            {8'h00}, /* 0x59ae */
            {8'h00}, /* 0x59ad */
            {8'h00}, /* 0x59ac */
            {8'h00}, /* 0x59ab */
            {8'h00}, /* 0x59aa */
            {8'h00}, /* 0x59a9 */
            {8'h00}, /* 0x59a8 */
            {8'h00}, /* 0x59a7 */
            {8'h00}, /* 0x59a6 */
            {8'h00}, /* 0x59a5 */
            {8'h00}, /* 0x59a4 */
            {8'h00}, /* 0x59a3 */
            {8'h00}, /* 0x59a2 */
            {8'h00}, /* 0x59a1 */
            {8'h00}, /* 0x59a0 */
            {8'h00}, /* 0x599f */
            {8'h00}, /* 0x599e */
            {8'h00}, /* 0x599d */
            {8'h00}, /* 0x599c */
            {8'h00}, /* 0x599b */
            {8'h00}, /* 0x599a */
            {8'h00}, /* 0x5999 */
            {8'h00}, /* 0x5998 */
            {8'h00}, /* 0x5997 */
            {8'h00}, /* 0x5996 */
            {8'h00}, /* 0x5995 */
            {8'h00}, /* 0x5994 */
            {8'h00}, /* 0x5993 */
            {8'h00}, /* 0x5992 */
            {8'h00}, /* 0x5991 */
            {8'h00}, /* 0x5990 */
            {8'h00}, /* 0x598f */
            {8'h00}, /* 0x598e */
            {8'h00}, /* 0x598d */
            {8'h00}, /* 0x598c */
            {8'h00}, /* 0x598b */
            {8'h00}, /* 0x598a */
            {8'h00}, /* 0x5989 */
            {8'h00}, /* 0x5988 */
            {8'h00}, /* 0x5987 */
            {8'h00}, /* 0x5986 */
            {8'h00}, /* 0x5985 */
            {8'h00}, /* 0x5984 */
            {8'h00}, /* 0x5983 */
            {8'h00}, /* 0x5982 */
            {8'h00}, /* 0x5981 */
            {8'h00}, /* 0x5980 */
            {8'h00}, /* 0x597f */
            {8'h00}, /* 0x597e */
            {8'h00}, /* 0x597d */
            {8'h00}, /* 0x597c */
            {8'h00}, /* 0x597b */
            {8'h00}, /* 0x597a */
            {8'h00}, /* 0x5979 */
            {8'h00}, /* 0x5978 */
            {8'h00}, /* 0x5977 */
            {8'h00}, /* 0x5976 */
            {8'h00}, /* 0x5975 */
            {8'h00}, /* 0x5974 */
            {8'h00}, /* 0x5973 */
            {8'h00}, /* 0x5972 */
            {8'h00}, /* 0x5971 */
            {8'h00}, /* 0x5970 */
            {8'h00}, /* 0x596f */
            {8'h00}, /* 0x596e */
            {8'h00}, /* 0x596d */
            {8'h00}, /* 0x596c */
            {8'h00}, /* 0x596b */
            {8'h00}, /* 0x596a */
            {8'h00}, /* 0x5969 */
            {8'h00}, /* 0x5968 */
            {8'h00}, /* 0x5967 */
            {8'h00}, /* 0x5966 */
            {8'h00}, /* 0x5965 */
            {8'h00}, /* 0x5964 */
            {8'h00}, /* 0x5963 */
            {8'h00}, /* 0x5962 */
            {8'h00}, /* 0x5961 */
            {8'h00}, /* 0x5960 */
            {8'h00}, /* 0x595f */
            {8'h00}, /* 0x595e */
            {8'h00}, /* 0x595d */
            {8'h00}, /* 0x595c */
            {8'h00}, /* 0x595b */
            {8'h00}, /* 0x595a */
            {8'h00}, /* 0x5959 */
            {8'h00}, /* 0x5958 */
            {8'h00}, /* 0x5957 */
            {8'h00}, /* 0x5956 */
            {8'h00}, /* 0x5955 */
            {8'h00}, /* 0x5954 */
            {8'h00}, /* 0x5953 */
            {8'h00}, /* 0x5952 */
            {8'h00}, /* 0x5951 */
            {8'h00}, /* 0x5950 */
            {8'h00}, /* 0x594f */
            {8'h00}, /* 0x594e */
            {8'h00}, /* 0x594d */
            {8'h00}, /* 0x594c */
            {8'h00}, /* 0x594b */
            {8'h00}, /* 0x594a */
            {8'h00}, /* 0x5949 */
            {8'h00}, /* 0x5948 */
            {8'h00}, /* 0x5947 */
            {8'h00}, /* 0x5946 */
            {8'h00}, /* 0x5945 */
            {8'h00}, /* 0x5944 */
            {8'h00}, /* 0x5943 */
            {8'h00}, /* 0x5942 */
            {8'h00}, /* 0x5941 */
            {8'h00}, /* 0x5940 */
            {8'h00}, /* 0x593f */
            {8'h00}, /* 0x593e */
            {8'h00}, /* 0x593d */
            {8'h00}, /* 0x593c */
            {8'h00}, /* 0x593b */
            {8'h00}, /* 0x593a */
            {8'h00}, /* 0x5939 */
            {8'h00}, /* 0x5938 */
            {8'h00}, /* 0x5937 */
            {8'h00}, /* 0x5936 */
            {8'h00}, /* 0x5935 */
            {8'h00}, /* 0x5934 */
            {8'h00}, /* 0x5933 */
            {8'h00}, /* 0x5932 */
            {8'h00}, /* 0x5931 */
            {8'h00}, /* 0x5930 */
            {8'h00}, /* 0x592f */
            {8'h00}, /* 0x592e */
            {8'h00}, /* 0x592d */
            {8'h00}, /* 0x592c */
            {8'h00}, /* 0x592b */
            {8'h00}, /* 0x592a */
            {8'h00}, /* 0x5929 */
            {8'h00}, /* 0x5928 */
            {8'h00}, /* 0x5927 */
            {8'h00}, /* 0x5926 */
            {8'h00}, /* 0x5925 */
            {8'h00}, /* 0x5924 */
            {8'h00}, /* 0x5923 */
            {8'h00}, /* 0x5922 */
            {8'h00}, /* 0x5921 */
            {8'h00}, /* 0x5920 */
            {8'h00}, /* 0x591f */
            {8'h00}, /* 0x591e */
            {8'h00}, /* 0x591d */
            {8'h00}, /* 0x591c */
            {8'h00}, /* 0x591b */
            {8'h00}, /* 0x591a */
            {8'h00}, /* 0x5919 */
            {8'h00}, /* 0x5918 */
            {8'h00}, /* 0x5917 */
            {8'h00}, /* 0x5916 */
            {8'h00}, /* 0x5915 */
            {8'h00}, /* 0x5914 */
            {8'h00}, /* 0x5913 */
            {8'h00}, /* 0x5912 */
            {8'h00}, /* 0x5911 */
            {8'h00}, /* 0x5910 */
            {8'h00}, /* 0x590f */
            {8'h00}, /* 0x590e */
            {8'h00}, /* 0x590d */
            {8'h00}, /* 0x590c */
            {8'h00}, /* 0x590b */
            {8'h00}, /* 0x590a */
            {8'h00}, /* 0x5909 */
            {8'h00}, /* 0x5908 */
            {8'h00}, /* 0x5907 */
            {8'h00}, /* 0x5906 */
            {8'h00}, /* 0x5905 */
            {8'h00}, /* 0x5904 */
            {8'h00}, /* 0x5903 */
            {8'h00}, /* 0x5902 */
            {8'h00}, /* 0x5901 */
            {8'h00}, /* 0x5900 */
            {8'h00}, /* 0x58ff */
            {8'h00}, /* 0x58fe */
            {8'h00}, /* 0x58fd */
            {8'h00}, /* 0x58fc */
            {8'h00}, /* 0x58fb */
            {8'h00}, /* 0x58fa */
            {8'h00}, /* 0x58f9 */
            {8'h00}, /* 0x58f8 */
            {8'h00}, /* 0x58f7 */
            {8'h00}, /* 0x58f6 */
            {8'h00}, /* 0x58f5 */
            {8'h00}, /* 0x58f4 */
            {8'h00}, /* 0x58f3 */
            {8'h00}, /* 0x58f2 */
            {8'h00}, /* 0x58f1 */
            {8'h00}, /* 0x58f0 */
            {8'h00}, /* 0x58ef */
            {8'h00}, /* 0x58ee */
            {8'h00}, /* 0x58ed */
            {8'h00}, /* 0x58ec */
            {8'h00}, /* 0x58eb */
            {8'h00}, /* 0x58ea */
            {8'h00}, /* 0x58e9 */
            {8'h00}, /* 0x58e8 */
            {8'h00}, /* 0x58e7 */
            {8'h00}, /* 0x58e6 */
            {8'h00}, /* 0x58e5 */
            {8'h00}, /* 0x58e4 */
            {8'h00}, /* 0x58e3 */
            {8'h00}, /* 0x58e2 */
            {8'h00}, /* 0x58e1 */
            {8'h00}, /* 0x58e0 */
            {8'h00}, /* 0x58df */
            {8'h00}, /* 0x58de */
            {8'h00}, /* 0x58dd */
            {8'h00}, /* 0x58dc */
            {8'h00}, /* 0x58db */
            {8'h00}, /* 0x58da */
            {8'h00}, /* 0x58d9 */
            {8'h00}, /* 0x58d8 */
            {8'h00}, /* 0x58d7 */
            {8'h00}, /* 0x58d6 */
            {8'h00}, /* 0x58d5 */
            {8'h00}, /* 0x58d4 */
            {8'h00}, /* 0x58d3 */
            {8'h00}, /* 0x58d2 */
            {8'h00}, /* 0x58d1 */
            {8'h00}, /* 0x58d0 */
            {8'h00}, /* 0x58cf */
            {8'h00}, /* 0x58ce */
            {8'h00}, /* 0x58cd */
            {8'h00}, /* 0x58cc */
            {8'h00}, /* 0x58cb */
            {8'h00}, /* 0x58ca */
            {8'h00}, /* 0x58c9 */
            {8'h00}, /* 0x58c8 */
            {8'h00}, /* 0x58c7 */
            {8'h00}, /* 0x58c6 */
            {8'h00}, /* 0x58c5 */
            {8'h00}, /* 0x58c4 */
            {8'h00}, /* 0x58c3 */
            {8'h00}, /* 0x58c2 */
            {8'h00}, /* 0x58c1 */
            {8'h00}, /* 0x58c0 */
            {8'h00}, /* 0x58bf */
            {8'h00}, /* 0x58be */
            {8'h00}, /* 0x58bd */
            {8'h00}, /* 0x58bc */
            {8'h00}, /* 0x58bb */
            {8'h00}, /* 0x58ba */
            {8'h00}, /* 0x58b9 */
            {8'h00}, /* 0x58b8 */
            {8'h00}, /* 0x58b7 */
            {8'h00}, /* 0x58b6 */
            {8'h00}, /* 0x58b5 */
            {8'h00}, /* 0x58b4 */
            {8'h00}, /* 0x58b3 */
            {8'h00}, /* 0x58b2 */
            {8'h00}, /* 0x58b1 */
            {8'h00}, /* 0x58b0 */
            {8'h00}, /* 0x58af */
            {8'h00}, /* 0x58ae */
            {8'h00}, /* 0x58ad */
            {8'h00}, /* 0x58ac */
            {8'h00}, /* 0x58ab */
            {8'h00}, /* 0x58aa */
            {8'h00}, /* 0x58a9 */
            {8'h00}, /* 0x58a8 */
            {8'h00}, /* 0x58a7 */
            {8'h00}, /* 0x58a6 */
            {8'h00}, /* 0x58a5 */
            {8'h00}, /* 0x58a4 */
            {8'h00}, /* 0x58a3 */
            {8'h00}, /* 0x58a2 */
            {8'h00}, /* 0x58a1 */
            {8'h00}, /* 0x58a0 */
            {8'h00}, /* 0x589f */
            {8'h00}, /* 0x589e */
            {8'h00}, /* 0x589d */
            {8'h00}, /* 0x589c */
            {8'h00}, /* 0x589b */
            {8'h00}, /* 0x589a */
            {8'h00}, /* 0x5899 */
            {8'h00}, /* 0x5898 */
            {8'h00}, /* 0x5897 */
            {8'h00}, /* 0x5896 */
            {8'h00}, /* 0x5895 */
            {8'h00}, /* 0x5894 */
            {8'h00}, /* 0x5893 */
            {8'h00}, /* 0x5892 */
            {8'h00}, /* 0x5891 */
            {8'h00}, /* 0x5890 */
            {8'h00}, /* 0x588f */
            {8'h00}, /* 0x588e */
            {8'h00}, /* 0x588d */
            {8'h00}, /* 0x588c */
            {8'h00}, /* 0x588b */
            {8'h00}, /* 0x588a */
            {8'h00}, /* 0x5889 */
            {8'h00}, /* 0x5888 */
            {8'h00}, /* 0x5887 */
            {8'h00}, /* 0x5886 */
            {8'h00}, /* 0x5885 */
            {8'h00}, /* 0x5884 */
            {8'h00}, /* 0x5883 */
            {8'h00}, /* 0x5882 */
            {8'h00}, /* 0x5881 */
            {8'h00}, /* 0x5880 */
            {8'h00}, /* 0x587f */
            {8'h00}, /* 0x587e */
            {8'h00}, /* 0x587d */
            {8'h00}, /* 0x587c */
            {8'h00}, /* 0x587b */
            {8'h00}, /* 0x587a */
            {8'h00}, /* 0x5879 */
            {8'h00}, /* 0x5878 */
            {8'h00}, /* 0x5877 */
            {8'h00}, /* 0x5876 */
            {8'h00}, /* 0x5875 */
            {8'h00}, /* 0x5874 */
            {8'h00}, /* 0x5873 */
            {8'h00}, /* 0x5872 */
            {8'h00}, /* 0x5871 */
            {8'h00}, /* 0x5870 */
            {8'h00}, /* 0x586f */
            {8'h00}, /* 0x586e */
            {8'h00}, /* 0x586d */
            {8'h00}, /* 0x586c */
            {8'h00}, /* 0x586b */
            {8'h00}, /* 0x586a */
            {8'h00}, /* 0x5869 */
            {8'h00}, /* 0x5868 */
            {8'h00}, /* 0x5867 */
            {8'h00}, /* 0x5866 */
            {8'h00}, /* 0x5865 */
            {8'h00}, /* 0x5864 */
            {8'h00}, /* 0x5863 */
            {8'h00}, /* 0x5862 */
            {8'h00}, /* 0x5861 */
            {8'h00}, /* 0x5860 */
            {8'h00}, /* 0x585f */
            {8'h00}, /* 0x585e */
            {8'h00}, /* 0x585d */
            {8'h00}, /* 0x585c */
            {8'h00}, /* 0x585b */
            {8'h00}, /* 0x585a */
            {8'h00}, /* 0x5859 */
            {8'h00}, /* 0x5858 */
            {8'h00}, /* 0x5857 */
            {8'h00}, /* 0x5856 */
            {8'h00}, /* 0x5855 */
            {8'h00}, /* 0x5854 */
            {8'h00}, /* 0x5853 */
            {8'h00}, /* 0x5852 */
            {8'h00}, /* 0x5851 */
            {8'h00}, /* 0x5850 */
            {8'h00}, /* 0x584f */
            {8'h00}, /* 0x584e */
            {8'h00}, /* 0x584d */
            {8'h00}, /* 0x584c */
            {8'h00}, /* 0x584b */
            {8'h00}, /* 0x584a */
            {8'h00}, /* 0x5849 */
            {8'h00}, /* 0x5848 */
            {8'h00}, /* 0x5847 */
            {8'h00}, /* 0x5846 */
            {8'h00}, /* 0x5845 */
            {8'h00}, /* 0x5844 */
            {8'h00}, /* 0x5843 */
            {8'h00}, /* 0x5842 */
            {8'h00}, /* 0x5841 */
            {8'h00}, /* 0x5840 */
            {8'h00}, /* 0x583f */
            {8'h00}, /* 0x583e */
            {8'h00}, /* 0x583d */
            {8'h00}, /* 0x583c */
            {8'h00}, /* 0x583b */
            {8'h00}, /* 0x583a */
            {8'h00}, /* 0x5839 */
            {8'h00}, /* 0x5838 */
            {8'h00}, /* 0x5837 */
            {8'h00}, /* 0x5836 */
            {8'h00}, /* 0x5835 */
            {8'h00}, /* 0x5834 */
            {8'h00}, /* 0x5833 */
            {8'h00}, /* 0x5832 */
            {8'h00}, /* 0x5831 */
            {8'h00}, /* 0x5830 */
            {8'h00}, /* 0x582f */
            {8'h00}, /* 0x582e */
            {8'h00}, /* 0x582d */
            {8'h00}, /* 0x582c */
            {8'h00}, /* 0x582b */
            {8'h00}, /* 0x582a */
            {8'h00}, /* 0x5829 */
            {8'h00}, /* 0x5828 */
            {8'h00}, /* 0x5827 */
            {8'h00}, /* 0x5826 */
            {8'h00}, /* 0x5825 */
            {8'h00}, /* 0x5824 */
            {8'h00}, /* 0x5823 */
            {8'h00}, /* 0x5822 */
            {8'h00}, /* 0x5821 */
            {8'h00}, /* 0x5820 */
            {8'h00}, /* 0x581f */
            {8'h00}, /* 0x581e */
            {8'h00}, /* 0x581d */
            {8'h00}, /* 0x581c */
            {8'h00}, /* 0x581b */
            {8'h00}, /* 0x581a */
            {8'h00}, /* 0x5819 */
            {8'h00}, /* 0x5818 */
            {8'h00}, /* 0x5817 */
            {8'h00}, /* 0x5816 */
            {8'h00}, /* 0x5815 */
            {8'h00}, /* 0x5814 */
            {8'h00}, /* 0x5813 */
            {8'h00}, /* 0x5812 */
            {8'h00}, /* 0x5811 */
            {8'h00}, /* 0x5810 */
            {8'h00}, /* 0x580f */
            {8'h00}, /* 0x580e */
            {8'h00}, /* 0x580d */
            {8'h00}, /* 0x580c */
            {8'h00}, /* 0x580b */
            {8'h00}, /* 0x580a */
            {8'h00}, /* 0x5809 */
            {8'h00}, /* 0x5808 */
            {8'h00}, /* 0x5807 */
            {8'h00}, /* 0x5806 */
            {8'h00}, /* 0x5805 */
            {8'h00}, /* 0x5804 */
            {8'h00}, /* 0x5803 */
            {8'h00}, /* 0x5802 */
            {8'h00}, /* 0x5801 */
            {8'h00}, /* 0x5800 */
            {8'h00}, /* 0x57ff */
            {8'h00}, /* 0x57fe */
            {8'h00}, /* 0x57fd */
            {8'h00}, /* 0x57fc */
            {8'h00}, /* 0x57fb */
            {8'h00}, /* 0x57fa */
            {8'h00}, /* 0x57f9 */
            {8'h00}, /* 0x57f8 */
            {8'h00}, /* 0x57f7 */
            {8'h00}, /* 0x57f6 */
            {8'h00}, /* 0x57f5 */
            {8'h00}, /* 0x57f4 */
            {8'h00}, /* 0x57f3 */
            {8'h00}, /* 0x57f2 */
            {8'h00}, /* 0x57f1 */
            {8'h00}, /* 0x57f0 */
            {8'h00}, /* 0x57ef */
            {8'h00}, /* 0x57ee */
            {8'h00}, /* 0x57ed */
            {8'h00}, /* 0x57ec */
            {8'h00}, /* 0x57eb */
            {8'h00}, /* 0x57ea */
            {8'h00}, /* 0x57e9 */
            {8'h00}, /* 0x57e8 */
            {8'h00}, /* 0x57e7 */
            {8'h00}, /* 0x57e6 */
            {8'h00}, /* 0x57e5 */
            {8'h00}, /* 0x57e4 */
            {8'h00}, /* 0x57e3 */
            {8'h00}, /* 0x57e2 */
            {8'h00}, /* 0x57e1 */
            {8'h00}, /* 0x57e0 */
            {8'h00}, /* 0x57df */
            {8'h00}, /* 0x57de */
            {8'h00}, /* 0x57dd */
            {8'h00}, /* 0x57dc */
            {8'h00}, /* 0x57db */
            {8'h00}, /* 0x57da */
            {8'h00}, /* 0x57d9 */
            {8'h00}, /* 0x57d8 */
            {8'h00}, /* 0x57d7 */
            {8'h00}, /* 0x57d6 */
            {8'h00}, /* 0x57d5 */
            {8'h00}, /* 0x57d4 */
            {8'h00}, /* 0x57d3 */
            {8'h00}, /* 0x57d2 */
            {8'h00}, /* 0x57d1 */
            {8'h00}, /* 0x57d0 */
            {8'h00}, /* 0x57cf */
            {8'h00}, /* 0x57ce */
            {8'h00}, /* 0x57cd */
            {8'h00}, /* 0x57cc */
            {8'h00}, /* 0x57cb */
            {8'h00}, /* 0x57ca */
            {8'h00}, /* 0x57c9 */
            {8'h00}, /* 0x57c8 */
            {8'h00}, /* 0x57c7 */
            {8'h00}, /* 0x57c6 */
            {8'h00}, /* 0x57c5 */
            {8'h00}, /* 0x57c4 */
            {8'h00}, /* 0x57c3 */
            {8'h00}, /* 0x57c2 */
            {8'h00}, /* 0x57c1 */
            {8'h00}, /* 0x57c0 */
            {8'h00}, /* 0x57bf */
            {8'h00}, /* 0x57be */
            {8'h00}, /* 0x57bd */
            {8'h00}, /* 0x57bc */
            {8'h00}, /* 0x57bb */
            {8'h00}, /* 0x57ba */
            {8'h00}, /* 0x57b9 */
            {8'h00}, /* 0x57b8 */
            {8'h00}, /* 0x57b7 */
            {8'h00}, /* 0x57b6 */
            {8'h00}, /* 0x57b5 */
            {8'h00}, /* 0x57b4 */
            {8'h00}, /* 0x57b3 */
            {8'h00}, /* 0x57b2 */
            {8'h00}, /* 0x57b1 */
            {8'h00}, /* 0x57b0 */
            {8'h00}, /* 0x57af */
            {8'h00}, /* 0x57ae */
            {8'h00}, /* 0x57ad */
            {8'h00}, /* 0x57ac */
            {8'h00}, /* 0x57ab */
            {8'h00}, /* 0x57aa */
            {8'h00}, /* 0x57a9 */
            {8'h00}, /* 0x57a8 */
            {8'h00}, /* 0x57a7 */
            {8'h00}, /* 0x57a6 */
            {8'h00}, /* 0x57a5 */
            {8'h00}, /* 0x57a4 */
            {8'h00}, /* 0x57a3 */
            {8'h00}, /* 0x57a2 */
            {8'h00}, /* 0x57a1 */
            {8'h00}, /* 0x57a0 */
            {8'h00}, /* 0x579f */
            {8'h00}, /* 0x579e */
            {8'h00}, /* 0x579d */
            {8'h00}, /* 0x579c */
            {8'h00}, /* 0x579b */
            {8'h00}, /* 0x579a */
            {8'h00}, /* 0x5799 */
            {8'h00}, /* 0x5798 */
            {8'h00}, /* 0x5797 */
            {8'h00}, /* 0x5796 */
            {8'h00}, /* 0x5795 */
            {8'h00}, /* 0x5794 */
            {8'h00}, /* 0x5793 */
            {8'h00}, /* 0x5792 */
            {8'h00}, /* 0x5791 */
            {8'h00}, /* 0x5790 */
            {8'h00}, /* 0x578f */
            {8'h00}, /* 0x578e */
            {8'h00}, /* 0x578d */
            {8'h00}, /* 0x578c */
            {8'h00}, /* 0x578b */
            {8'h00}, /* 0x578a */
            {8'h00}, /* 0x5789 */
            {8'h00}, /* 0x5788 */
            {8'h00}, /* 0x5787 */
            {8'h00}, /* 0x5786 */
            {8'h00}, /* 0x5785 */
            {8'h00}, /* 0x5784 */
            {8'h00}, /* 0x5783 */
            {8'h00}, /* 0x5782 */
            {8'h00}, /* 0x5781 */
            {8'h00}, /* 0x5780 */
            {8'h00}, /* 0x577f */
            {8'h00}, /* 0x577e */
            {8'h00}, /* 0x577d */
            {8'h00}, /* 0x577c */
            {8'h00}, /* 0x577b */
            {8'h00}, /* 0x577a */
            {8'h00}, /* 0x5779 */
            {8'h00}, /* 0x5778 */
            {8'h00}, /* 0x5777 */
            {8'h00}, /* 0x5776 */
            {8'h00}, /* 0x5775 */
            {8'h00}, /* 0x5774 */
            {8'h00}, /* 0x5773 */
            {8'h00}, /* 0x5772 */
            {8'h00}, /* 0x5771 */
            {8'h00}, /* 0x5770 */
            {8'h00}, /* 0x576f */
            {8'h00}, /* 0x576e */
            {8'h00}, /* 0x576d */
            {8'h00}, /* 0x576c */
            {8'h00}, /* 0x576b */
            {8'h00}, /* 0x576a */
            {8'h00}, /* 0x5769 */
            {8'h00}, /* 0x5768 */
            {8'h00}, /* 0x5767 */
            {8'h00}, /* 0x5766 */
            {8'h00}, /* 0x5765 */
            {8'h00}, /* 0x5764 */
            {8'h00}, /* 0x5763 */
            {8'h00}, /* 0x5762 */
            {8'h00}, /* 0x5761 */
            {8'h00}, /* 0x5760 */
            {8'h00}, /* 0x575f */
            {8'h00}, /* 0x575e */
            {8'h00}, /* 0x575d */
            {8'h00}, /* 0x575c */
            {8'h00}, /* 0x575b */
            {8'h00}, /* 0x575a */
            {8'h00}, /* 0x5759 */
            {8'h00}, /* 0x5758 */
            {8'h00}, /* 0x5757 */
            {8'h00}, /* 0x5756 */
            {8'h00}, /* 0x5755 */
            {8'h00}, /* 0x5754 */
            {8'h00}, /* 0x5753 */
            {8'h00}, /* 0x5752 */
            {8'h00}, /* 0x5751 */
            {8'h00}, /* 0x5750 */
            {8'h00}, /* 0x574f */
            {8'h00}, /* 0x574e */
            {8'h00}, /* 0x574d */
            {8'h00}, /* 0x574c */
            {8'h00}, /* 0x574b */
            {8'h00}, /* 0x574a */
            {8'h00}, /* 0x5749 */
            {8'h00}, /* 0x5748 */
            {8'h00}, /* 0x5747 */
            {8'h00}, /* 0x5746 */
            {8'h00}, /* 0x5745 */
            {8'h00}, /* 0x5744 */
            {8'h00}, /* 0x5743 */
            {8'h00}, /* 0x5742 */
            {8'h00}, /* 0x5741 */
            {8'h00}, /* 0x5740 */
            {8'h00}, /* 0x573f */
            {8'h00}, /* 0x573e */
            {8'h00}, /* 0x573d */
            {8'h00}, /* 0x573c */
            {8'h00}, /* 0x573b */
            {8'h00}, /* 0x573a */
            {8'h00}, /* 0x5739 */
            {8'h00}, /* 0x5738 */
            {8'h00}, /* 0x5737 */
            {8'h00}, /* 0x5736 */
            {8'h00}, /* 0x5735 */
            {8'h00}, /* 0x5734 */
            {8'h00}, /* 0x5733 */
            {8'h00}, /* 0x5732 */
            {8'h00}, /* 0x5731 */
            {8'h00}, /* 0x5730 */
            {8'h00}, /* 0x572f */
            {8'h00}, /* 0x572e */
            {8'h00}, /* 0x572d */
            {8'h00}, /* 0x572c */
            {8'h00}, /* 0x572b */
            {8'h00}, /* 0x572a */
            {8'h00}, /* 0x5729 */
            {8'h00}, /* 0x5728 */
            {8'h00}, /* 0x5727 */
            {8'h00}, /* 0x5726 */
            {8'h00}, /* 0x5725 */
            {8'h00}, /* 0x5724 */
            {8'h00}, /* 0x5723 */
            {8'h00}, /* 0x5722 */
            {8'h00}, /* 0x5721 */
            {8'h00}, /* 0x5720 */
            {8'h00}, /* 0x571f */
            {8'h00}, /* 0x571e */
            {8'h00}, /* 0x571d */
            {8'h00}, /* 0x571c */
            {8'h00}, /* 0x571b */
            {8'h00}, /* 0x571a */
            {8'h00}, /* 0x5719 */
            {8'h00}, /* 0x5718 */
            {8'h00}, /* 0x5717 */
            {8'h00}, /* 0x5716 */
            {8'h00}, /* 0x5715 */
            {8'h00}, /* 0x5714 */
            {8'h00}, /* 0x5713 */
            {8'h00}, /* 0x5712 */
            {8'h00}, /* 0x5711 */
            {8'h00}, /* 0x5710 */
            {8'h00}, /* 0x570f */
            {8'h00}, /* 0x570e */
            {8'h00}, /* 0x570d */
            {8'h00}, /* 0x570c */
            {8'h00}, /* 0x570b */
            {8'h00}, /* 0x570a */
            {8'h00}, /* 0x5709 */
            {8'h00}, /* 0x5708 */
            {8'h00}, /* 0x5707 */
            {8'h00}, /* 0x5706 */
            {8'h00}, /* 0x5705 */
            {8'h00}, /* 0x5704 */
            {8'h00}, /* 0x5703 */
            {8'h00}, /* 0x5702 */
            {8'h00}, /* 0x5701 */
            {8'h00}, /* 0x5700 */
            {8'h00}, /* 0x56ff */
            {8'h00}, /* 0x56fe */
            {8'h00}, /* 0x56fd */
            {8'h00}, /* 0x56fc */
            {8'h00}, /* 0x56fb */
            {8'h00}, /* 0x56fa */
            {8'h00}, /* 0x56f9 */
            {8'h00}, /* 0x56f8 */
            {8'h00}, /* 0x56f7 */
            {8'h00}, /* 0x56f6 */
            {8'h00}, /* 0x56f5 */
            {8'h00}, /* 0x56f4 */
            {8'h00}, /* 0x56f3 */
            {8'h00}, /* 0x56f2 */
            {8'h00}, /* 0x56f1 */
            {8'h00}, /* 0x56f0 */
            {8'h00}, /* 0x56ef */
            {8'h00}, /* 0x56ee */
            {8'h00}, /* 0x56ed */
            {8'h00}, /* 0x56ec */
            {8'h00}, /* 0x56eb */
            {8'h00}, /* 0x56ea */
            {8'h00}, /* 0x56e9 */
            {8'h00}, /* 0x56e8 */
            {8'h00}, /* 0x56e7 */
            {8'h00}, /* 0x56e6 */
            {8'h00}, /* 0x56e5 */
            {8'h00}, /* 0x56e4 */
            {8'h00}, /* 0x56e3 */
            {8'h00}, /* 0x56e2 */
            {8'h00}, /* 0x56e1 */
            {8'h00}, /* 0x56e0 */
            {8'h00}, /* 0x56df */
            {8'h00}, /* 0x56de */
            {8'h00}, /* 0x56dd */
            {8'h00}, /* 0x56dc */
            {8'h00}, /* 0x56db */
            {8'h00}, /* 0x56da */
            {8'h00}, /* 0x56d9 */
            {8'h00}, /* 0x56d8 */
            {8'h00}, /* 0x56d7 */
            {8'h00}, /* 0x56d6 */
            {8'h00}, /* 0x56d5 */
            {8'h00}, /* 0x56d4 */
            {8'h00}, /* 0x56d3 */
            {8'h00}, /* 0x56d2 */
            {8'h00}, /* 0x56d1 */
            {8'h00}, /* 0x56d0 */
            {8'h00}, /* 0x56cf */
            {8'h00}, /* 0x56ce */
            {8'h00}, /* 0x56cd */
            {8'h00}, /* 0x56cc */
            {8'h00}, /* 0x56cb */
            {8'h00}, /* 0x56ca */
            {8'h00}, /* 0x56c9 */
            {8'h00}, /* 0x56c8 */
            {8'h00}, /* 0x56c7 */
            {8'h00}, /* 0x56c6 */
            {8'h00}, /* 0x56c5 */
            {8'h00}, /* 0x56c4 */
            {8'h00}, /* 0x56c3 */
            {8'h00}, /* 0x56c2 */
            {8'h00}, /* 0x56c1 */
            {8'h00}, /* 0x56c0 */
            {8'h00}, /* 0x56bf */
            {8'h00}, /* 0x56be */
            {8'h00}, /* 0x56bd */
            {8'h00}, /* 0x56bc */
            {8'h00}, /* 0x56bb */
            {8'h00}, /* 0x56ba */
            {8'h00}, /* 0x56b9 */
            {8'h00}, /* 0x56b8 */
            {8'h00}, /* 0x56b7 */
            {8'h00}, /* 0x56b6 */
            {8'h00}, /* 0x56b5 */
            {8'h00}, /* 0x56b4 */
            {8'h00}, /* 0x56b3 */
            {8'h00}, /* 0x56b2 */
            {8'h00}, /* 0x56b1 */
            {8'h00}, /* 0x56b0 */
            {8'h00}, /* 0x56af */
            {8'h00}, /* 0x56ae */
            {8'h00}, /* 0x56ad */
            {8'h00}, /* 0x56ac */
            {8'h00}, /* 0x56ab */
            {8'h00}, /* 0x56aa */
            {8'h00}, /* 0x56a9 */
            {8'h00}, /* 0x56a8 */
            {8'h00}, /* 0x56a7 */
            {8'h00}, /* 0x56a6 */
            {8'h00}, /* 0x56a5 */
            {8'h00}, /* 0x56a4 */
            {8'h00}, /* 0x56a3 */
            {8'h00}, /* 0x56a2 */
            {8'h00}, /* 0x56a1 */
            {8'h00}, /* 0x56a0 */
            {8'h00}, /* 0x569f */
            {8'h00}, /* 0x569e */
            {8'h00}, /* 0x569d */
            {8'h00}, /* 0x569c */
            {8'h00}, /* 0x569b */
            {8'h00}, /* 0x569a */
            {8'h00}, /* 0x5699 */
            {8'h00}, /* 0x5698 */
            {8'h00}, /* 0x5697 */
            {8'h00}, /* 0x5696 */
            {8'h00}, /* 0x5695 */
            {8'h00}, /* 0x5694 */
            {8'h00}, /* 0x5693 */
            {8'h00}, /* 0x5692 */
            {8'h00}, /* 0x5691 */
            {8'h00}, /* 0x5690 */
            {8'h00}, /* 0x568f */
            {8'h00}, /* 0x568e */
            {8'h00}, /* 0x568d */
            {8'h00}, /* 0x568c */
            {8'h00}, /* 0x568b */
            {8'h00}, /* 0x568a */
            {8'h00}, /* 0x5689 */
            {8'h00}, /* 0x5688 */
            {8'h00}, /* 0x5687 */
            {8'h00}, /* 0x5686 */
            {8'h00}, /* 0x5685 */
            {8'h00}, /* 0x5684 */
            {8'h00}, /* 0x5683 */
            {8'h00}, /* 0x5682 */
            {8'h00}, /* 0x5681 */
            {8'h00}, /* 0x5680 */
            {8'h00}, /* 0x567f */
            {8'h00}, /* 0x567e */
            {8'h00}, /* 0x567d */
            {8'h00}, /* 0x567c */
            {8'h00}, /* 0x567b */
            {8'h00}, /* 0x567a */
            {8'h00}, /* 0x5679 */
            {8'h00}, /* 0x5678 */
            {8'h00}, /* 0x5677 */
            {8'h00}, /* 0x5676 */
            {8'h00}, /* 0x5675 */
            {8'h00}, /* 0x5674 */
            {8'h00}, /* 0x5673 */
            {8'h00}, /* 0x5672 */
            {8'h00}, /* 0x5671 */
            {8'h00}, /* 0x5670 */
            {8'h00}, /* 0x566f */
            {8'h00}, /* 0x566e */
            {8'h00}, /* 0x566d */
            {8'h00}, /* 0x566c */
            {8'h00}, /* 0x566b */
            {8'h00}, /* 0x566a */
            {8'h00}, /* 0x5669 */
            {8'h00}, /* 0x5668 */
            {8'h00}, /* 0x5667 */
            {8'h00}, /* 0x5666 */
            {8'h00}, /* 0x5665 */
            {8'h00}, /* 0x5664 */
            {8'h00}, /* 0x5663 */
            {8'h00}, /* 0x5662 */
            {8'h00}, /* 0x5661 */
            {8'h00}, /* 0x5660 */
            {8'h00}, /* 0x565f */
            {8'h00}, /* 0x565e */
            {8'h00}, /* 0x565d */
            {8'h00}, /* 0x565c */
            {8'h00}, /* 0x565b */
            {8'h00}, /* 0x565a */
            {8'h00}, /* 0x5659 */
            {8'h00}, /* 0x5658 */
            {8'h00}, /* 0x5657 */
            {8'h00}, /* 0x5656 */
            {8'h00}, /* 0x5655 */
            {8'h00}, /* 0x5654 */
            {8'h00}, /* 0x5653 */
            {8'h00}, /* 0x5652 */
            {8'h00}, /* 0x5651 */
            {8'h00}, /* 0x5650 */
            {8'h00}, /* 0x564f */
            {8'h00}, /* 0x564e */
            {8'h00}, /* 0x564d */
            {8'h00}, /* 0x564c */
            {8'h00}, /* 0x564b */
            {8'h00}, /* 0x564a */
            {8'h00}, /* 0x5649 */
            {8'h00}, /* 0x5648 */
            {8'h00}, /* 0x5647 */
            {8'h00}, /* 0x5646 */
            {8'h00}, /* 0x5645 */
            {8'h00}, /* 0x5644 */
            {8'h00}, /* 0x5643 */
            {8'h00}, /* 0x5642 */
            {8'h00}, /* 0x5641 */
            {8'h00}, /* 0x5640 */
            {8'h00}, /* 0x563f */
            {8'h00}, /* 0x563e */
            {8'h00}, /* 0x563d */
            {8'h00}, /* 0x563c */
            {8'h00}, /* 0x563b */
            {8'h00}, /* 0x563a */
            {8'h00}, /* 0x5639 */
            {8'h00}, /* 0x5638 */
            {8'h00}, /* 0x5637 */
            {8'h00}, /* 0x5636 */
            {8'h00}, /* 0x5635 */
            {8'h00}, /* 0x5634 */
            {8'h00}, /* 0x5633 */
            {8'h00}, /* 0x5632 */
            {8'h00}, /* 0x5631 */
            {8'h00}, /* 0x5630 */
            {8'h00}, /* 0x562f */
            {8'h00}, /* 0x562e */
            {8'h00}, /* 0x562d */
            {8'h00}, /* 0x562c */
            {8'h00}, /* 0x562b */
            {8'h00}, /* 0x562a */
            {8'h00}, /* 0x5629 */
            {8'h00}, /* 0x5628 */
            {8'h00}, /* 0x5627 */
            {8'h00}, /* 0x5626 */
            {8'h00}, /* 0x5625 */
            {8'h00}, /* 0x5624 */
            {8'h00}, /* 0x5623 */
            {8'h00}, /* 0x5622 */
            {8'h00}, /* 0x5621 */
            {8'h00}, /* 0x5620 */
            {8'h00}, /* 0x561f */
            {8'h00}, /* 0x561e */
            {8'h00}, /* 0x561d */
            {8'h00}, /* 0x561c */
            {8'h00}, /* 0x561b */
            {8'h00}, /* 0x561a */
            {8'h00}, /* 0x5619 */
            {8'h00}, /* 0x5618 */
            {8'h00}, /* 0x5617 */
            {8'h00}, /* 0x5616 */
            {8'h00}, /* 0x5615 */
            {8'h00}, /* 0x5614 */
            {8'h00}, /* 0x5613 */
            {8'h00}, /* 0x5612 */
            {8'h00}, /* 0x5611 */
            {8'h00}, /* 0x5610 */
            {8'h00}, /* 0x560f */
            {8'h00}, /* 0x560e */
            {8'h00}, /* 0x560d */
            {8'h00}, /* 0x560c */
            {8'h00}, /* 0x560b */
            {8'h00}, /* 0x560a */
            {8'h00}, /* 0x5609 */
            {8'h00}, /* 0x5608 */
            {8'h00}, /* 0x5607 */
            {8'h00}, /* 0x5606 */
            {8'h00}, /* 0x5605 */
            {8'h00}, /* 0x5604 */
            {8'h00}, /* 0x5603 */
            {8'h00}, /* 0x5602 */
            {8'h00}, /* 0x5601 */
            {8'h00}, /* 0x5600 */
            {8'h00}, /* 0x55ff */
            {8'h00}, /* 0x55fe */
            {8'h00}, /* 0x55fd */
            {8'h00}, /* 0x55fc */
            {8'h00}, /* 0x55fb */
            {8'h00}, /* 0x55fa */
            {8'h00}, /* 0x55f9 */
            {8'h00}, /* 0x55f8 */
            {8'h00}, /* 0x55f7 */
            {8'h00}, /* 0x55f6 */
            {8'h00}, /* 0x55f5 */
            {8'h00}, /* 0x55f4 */
            {8'h00}, /* 0x55f3 */
            {8'h00}, /* 0x55f2 */
            {8'h00}, /* 0x55f1 */
            {8'h00}, /* 0x55f0 */
            {8'h00}, /* 0x55ef */
            {8'h00}, /* 0x55ee */
            {8'h00}, /* 0x55ed */
            {8'h00}, /* 0x55ec */
            {8'h00}, /* 0x55eb */
            {8'h00}, /* 0x55ea */
            {8'h00}, /* 0x55e9 */
            {8'h00}, /* 0x55e8 */
            {8'h00}, /* 0x55e7 */
            {8'h00}, /* 0x55e6 */
            {8'h00}, /* 0x55e5 */
            {8'h00}, /* 0x55e4 */
            {8'h00}, /* 0x55e3 */
            {8'h00}, /* 0x55e2 */
            {8'h00}, /* 0x55e1 */
            {8'h00}, /* 0x55e0 */
            {8'h00}, /* 0x55df */
            {8'h00}, /* 0x55de */
            {8'h00}, /* 0x55dd */
            {8'h00}, /* 0x55dc */
            {8'h00}, /* 0x55db */
            {8'h00}, /* 0x55da */
            {8'h00}, /* 0x55d9 */
            {8'h00}, /* 0x55d8 */
            {8'h00}, /* 0x55d7 */
            {8'h00}, /* 0x55d6 */
            {8'h00}, /* 0x55d5 */
            {8'h00}, /* 0x55d4 */
            {8'h00}, /* 0x55d3 */
            {8'h00}, /* 0x55d2 */
            {8'h00}, /* 0x55d1 */
            {8'h00}, /* 0x55d0 */
            {8'h00}, /* 0x55cf */
            {8'h00}, /* 0x55ce */
            {8'h00}, /* 0x55cd */
            {8'h00}, /* 0x55cc */
            {8'h00}, /* 0x55cb */
            {8'h00}, /* 0x55ca */
            {8'h00}, /* 0x55c9 */
            {8'h00}, /* 0x55c8 */
            {8'h00}, /* 0x55c7 */
            {8'h00}, /* 0x55c6 */
            {8'h00}, /* 0x55c5 */
            {8'h00}, /* 0x55c4 */
            {8'h00}, /* 0x55c3 */
            {8'h00}, /* 0x55c2 */
            {8'h00}, /* 0x55c1 */
            {8'h00}, /* 0x55c0 */
            {8'h00}, /* 0x55bf */
            {8'h00}, /* 0x55be */
            {8'h00}, /* 0x55bd */
            {8'h00}, /* 0x55bc */
            {8'h00}, /* 0x55bb */
            {8'h00}, /* 0x55ba */
            {8'h00}, /* 0x55b9 */
            {8'h00}, /* 0x55b8 */
            {8'h00}, /* 0x55b7 */
            {8'h00}, /* 0x55b6 */
            {8'h00}, /* 0x55b5 */
            {8'h00}, /* 0x55b4 */
            {8'h00}, /* 0x55b3 */
            {8'h00}, /* 0x55b2 */
            {8'h00}, /* 0x55b1 */
            {8'h00}, /* 0x55b0 */
            {8'h00}, /* 0x55af */
            {8'h00}, /* 0x55ae */
            {8'h00}, /* 0x55ad */
            {8'h00}, /* 0x55ac */
            {8'h00}, /* 0x55ab */
            {8'h00}, /* 0x55aa */
            {8'h00}, /* 0x55a9 */
            {8'h00}, /* 0x55a8 */
            {8'h00}, /* 0x55a7 */
            {8'h00}, /* 0x55a6 */
            {8'h00}, /* 0x55a5 */
            {8'h00}, /* 0x55a4 */
            {8'h00}, /* 0x55a3 */
            {8'h00}, /* 0x55a2 */
            {8'h00}, /* 0x55a1 */
            {8'h00}, /* 0x55a0 */
            {8'h00}, /* 0x559f */
            {8'h00}, /* 0x559e */
            {8'h00}, /* 0x559d */
            {8'h00}, /* 0x559c */
            {8'h00}, /* 0x559b */
            {8'h00}, /* 0x559a */
            {8'h00}, /* 0x5599 */
            {8'h00}, /* 0x5598 */
            {8'h00}, /* 0x5597 */
            {8'h00}, /* 0x5596 */
            {8'h00}, /* 0x5595 */
            {8'h00}, /* 0x5594 */
            {8'h00}, /* 0x5593 */
            {8'h00}, /* 0x5592 */
            {8'h00}, /* 0x5591 */
            {8'h00}, /* 0x5590 */
            {8'h00}, /* 0x558f */
            {8'h00}, /* 0x558e */
            {8'h00}, /* 0x558d */
            {8'h00}, /* 0x558c */
            {8'h00}, /* 0x558b */
            {8'h00}, /* 0x558a */
            {8'h00}, /* 0x5589 */
            {8'h00}, /* 0x5588 */
            {8'h00}, /* 0x5587 */
            {8'h00}, /* 0x5586 */
            {8'h00}, /* 0x5585 */
            {8'h00}, /* 0x5584 */
            {8'h00}, /* 0x5583 */
            {8'h00}, /* 0x5582 */
            {8'h00}, /* 0x5581 */
            {8'h00}, /* 0x5580 */
            {8'h00}, /* 0x557f */
            {8'h00}, /* 0x557e */
            {8'h00}, /* 0x557d */
            {8'h00}, /* 0x557c */
            {8'h00}, /* 0x557b */
            {8'h00}, /* 0x557a */
            {8'h00}, /* 0x5579 */
            {8'h00}, /* 0x5578 */
            {8'h00}, /* 0x5577 */
            {8'h00}, /* 0x5576 */
            {8'h00}, /* 0x5575 */
            {8'h00}, /* 0x5574 */
            {8'h00}, /* 0x5573 */
            {8'h00}, /* 0x5572 */
            {8'h00}, /* 0x5571 */
            {8'h00}, /* 0x5570 */
            {8'h00}, /* 0x556f */
            {8'h00}, /* 0x556e */
            {8'h00}, /* 0x556d */
            {8'h00}, /* 0x556c */
            {8'h00}, /* 0x556b */
            {8'h00}, /* 0x556a */
            {8'h00}, /* 0x5569 */
            {8'h00}, /* 0x5568 */
            {8'h00}, /* 0x5567 */
            {8'h00}, /* 0x5566 */
            {8'h00}, /* 0x5565 */
            {8'h00}, /* 0x5564 */
            {8'h00}, /* 0x5563 */
            {8'h00}, /* 0x5562 */
            {8'h00}, /* 0x5561 */
            {8'h00}, /* 0x5560 */
            {8'h00}, /* 0x555f */
            {8'h00}, /* 0x555e */
            {8'h00}, /* 0x555d */
            {8'h00}, /* 0x555c */
            {8'h00}, /* 0x555b */
            {8'h00}, /* 0x555a */
            {8'h00}, /* 0x5559 */
            {8'h00}, /* 0x5558 */
            {8'h00}, /* 0x5557 */
            {8'h00}, /* 0x5556 */
            {8'h00}, /* 0x5555 */
            {8'h00}, /* 0x5554 */
            {8'h00}, /* 0x5553 */
            {8'h00}, /* 0x5552 */
            {8'h00}, /* 0x5551 */
            {8'h00}, /* 0x5550 */
            {8'h00}, /* 0x554f */
            {8'h00}, /* 0x554e */
            {8'h00}, /* 0x554d */
            {8'h00}, /* 0x554c */
            {8'h00}, /* 0x554b */
            {8'h00}, /* 0x554a */
            {8'h00}, /* 0x5549 */
            {8'h00}, /* 0x5548 */
            {8'h00}, /* 0x5547 */
            {8'h00}, /* 0x5546 */
            {8'h00}, /* 0x5545 */
            {8'h00}, /* 0x5544 */
            {8'h00}, /* 0x5543 */
            {8'h00}, /* 0x5542 */
            {8'h00}, /* 0x5541 */
            {8'h00}, /* 0x5540 */
            {8'h00}, /* 0x553f */
            {8'h00}, /* 0x553e */
            {8'h00}, /* 0x553d */
            {8'h00}, /* 0x553c */
            {8'h00}, /* 0x553b */
            {8'h00}, /* 0x553a */
            {8'h00}, /* 0x5539 */
            {8'h00}, /* 0x5538 */
            {8'h00}, /* 0x5537 */
            {8'h00}, /* 0x5536 */
            {8'h00}, /* 0x5535 */
            {8'h00}, /* 0x5534 */
            {8'h00}, /* 0x5533 */
            {8'h00}, /* 0x5532 */
            {8'h00}, /* 0x5531 */
            {8'h00}, /* 0x5530 */
            {8'h00}, /* 0x552f */
            {8'h00}, /* 0x552e */
            {8'h00}, /* 0x552d */
            {8'h00}, /* 0x552c */
            {8'h00}, /* 0x552b */
            {8'h00}, /* 0x552a */
            {8'h00}, /* 0x5529 */
            {8'h00}, /* 0x5528 */
            {8'h00}, /* 0x5527 */
            {8'h00}, /* 0x5526 */
            {8'h00}, /* 0x5525 */
            {8'h00}, /* 0x5524 */
            {8'h00}, /* 0x5523 */
            {8'h00}, /* 0x5522 */
            {8'h00}, /* 0x5521 */
            {8'h00}, /* 0x5520 */
            {8'h00}, /* 0x551f */
            {8'h00}, /* 0x551e */
            {8'h00}, /* 0x551d */
            {8'h00}, /* 0x551c */
            {8'h00}, /* 0x551b */
            {8'h00}, /* 0x551a */
            {8'h00}, /* 0x5519 */
            {8'h00}, /* 0x5518 */
            {8'h00}, /* 0x5517 */
            {8'h00}, /* 0x5516 */
            {8'h00}, /* 0x5515 */
            {8'h00}, /* 0x5514 */
            {8'h00}, /* 0x5513 */
            {8'h00}, /* 0x5512 */
            {8'h00}, /* 0x5511 */
            {8'h00}, /* 0x5510 */
            {8'h00}, /* 0x550f */
            {8'h00}, /* 0x550e */
            {8'h00}, /* 0x550d */
            {8'h00}, /* 0x550c */
            {8'h00}, /* 0x550b */
            {8'h00}, /* 0x550a */
            {8'h00}, /* 0x5509 */
            {8'h00}, /* 0x5508 */
            {8'h00}, /* 0x5507 */
            {8'h00}, /* 0x5506 */
            {8'h00}, /* 0x5505 */
            {8'h00}, /* 0x5504 */
            {8'h00}, /* 0x5503 */
            {8'h00}, /* 0x5502 */
            {8'h00}, /* 0x5501 */
            {8'h00}, /* 0x5500 */
            {8'h00}, /* 0x54ff */
            {8'h00}, /* 0x54fe */
            {8'h00}, /* 0x54fd */
            {8'h00}, /* 0x54fc */
            {8'h00}, /* 0x54fb */
            {8'h00}, /* 0x54fa */
            {8'h00}, /* 0x54f9 */
            {8'h00}, /* 0x54f8 */
            {8'h00}, /* 0x54f7 */
            {8'h00}, /* 0x54f6 */
            {8'h00}, /* 0x54f5 */
            {8'h00}, /* 0x54f4 */
            {8'h00}, /* 0x54f3 */
            {8'h00}, /* 0x54f2 */
            {8'h00}, /* 0x54f1 */
            {8'h00}, /* 0x54f0 */
            {8'h00}, /* 0x54ef */
            {8'h00}, /* 0x54ee */
            {8'h00}, /* 0x54ed */
            {8'h00}, /* 0x54ec */
            {8'h00}, /* 0x54eb */
            {8'h00}, /* 0x54ea */
            {8'h00}, /* 0x54e9 */
            {8'h00}, /* 0x54e8 */
            {8'h00}, /* 0x54e7 */
            {8'h00}, /* 0x54e6 */
            {8'h00}, /* 0x54e5 */
            {8'h00}, /* 0x54e4 */
            {8'h00}, /* 0x54e3 */
            {8'h00}, /* 0x54e2 */
            {8'h00}, /* 0x54e1 */
            {8'h00}, /* 0x54e0 */
            {8'h00}, /* 0x54df */
            {8'h00}, /* 0x54de */
            {8'h00}, /* 0x54dd */
            {8'h00}, /* 0x54dc */
            {8'h00}, /* 0x54db */
            {8'h00}, /* 0x54da */
            {8'h00}, /* 0x54d9 */
            {8'h00}, /* 0x54d8 */
            {8'h00}, /* 0x54d7 */
            {8'h00}, /* 0x54d6 */
            {8'h00}, /* 0x54d5 */
            {8'h00}, /* 0x54d4 */
            {8'h00}, /* 0x54d3 */
            {8'h00}, /* 0x54d2 */
            {8'h00}, /* 0x54d1 */
            {8'h00}, /* 0x54d0 */
            {8'h00}, /* 0x54cf */
            {8'h00}, /* 0x54ce */
            {8'h00}, /* 0x54cd */
            {8'h00}, /* 0x54cc */
            {8'h00}, /* 0x54cb */
            {8'h00}, /* 0x54ca */
            {8'h00}, /* 0x54c9 */
            {8'h00}, /* 0x54c8 */
            {8'h00}, /* 0x54c7 */
            {8'h00}, /* 0x54c6 */
            {8'h00}, /* 0x54c5 */
            {8'h00}, /* 0x54c4 */
            {8'h00}, /* 0x54c3 */
            {8'h00}, /* 0x54c2 */
            {8'h00}, /* 0x54c1 */
            {8'h00}, /* 0x54c0 */
            {8'h00}, /* 0x54bf */
            {8'h00}, /* 0x54be */
            {8'h00}, /* 0x54bd */
            {8'h00}, /* 0x54bc */
            {8'h00}, /* 0x54bb */
            {8'h00}, /* 0x54ba */
            {8'h00}, /* 0x54b9 */
            {8'h00}, /* 0x54b8 */
            {8'h00}, /* 0x54b7 */
            {8'h00}, /* 0x54b6 */
            {8'h00}, /* 0x54b5 */
            {8'h00}, /* 0x54b4 */
            {8'h00}, /* 0x54b3 */
            {8'h00}, /* 0x54b2 */
            {8'h00}, /* 0x54b1 */
            {8'h00}, /* 0x54b0 */
            {8'h00}, /* 0x54af */
            {8'h00}, /* 0x54ae */
            {8'h00}, /* 0x54ad */
            {8'h00}, /* 0x54ac */
            {8'h00}, /* 0x54ab */
            {8'h00}, /* 0x54aa */
            {8'h00}, /* 0x54a9 */
            {8'h00}, /* 0x54a8 */
            {8'h00}, /* 0x54a7 */
            {8'h00}, /* 0x54a6 */
            {8'h00}, /* 0x54a5 */
            {8'h00}, /* 0x54a4 */
            {8'h00}, /* 0x54a3 */
            {8'h00}, /* 0x54a2 */
            {8'h00}, /* 0x54a1 */
            {8'h00}, /* 0x54a0 */
            {8'h00}, /* 0x549f */
            {8'h00}, /* 0x549e */
            {8'h00}, /* 0x549d */
            {8'h00}, /* 0x549c */
            {8'h00}, /* 0x549b */
            {8'h00}, /* 0x549a */
            {8'h00}, /* 0x5499 */
            {8'h00}, /* 0x5498 */
            {8'h00}, /* 0x5497 */
            {8'h00}, /* 0x5496 */
            {8'h00}, /* 0x5495 */
            {8'h00}, /* 0x5494 */
            {8'h00}, /* 0x5493 */
            {8'h00}, /* 0x5492 */
            {8'h00}, /* 0x5491 */
            {8'h00}, /* 0x5490 */
            {8'h00}, /* 0x548f */
            {8'h00}, /* 0x548e */
            {8'h00}, /* 0x548d */
            {8'h00}, /* 0x548c */
            {8'h00}, /* 0x548b */
            {8'h00}, /* 0x548a */
            {8'h00}, /* 0x5489 */
            {8'h00}, /* 0x5488 */
            {8'h00}, /* 0x5487 */
            {8'h00}, /* 0x5486 */
            {8'h00}, /* 0x5485 */
            {8'h00}, /* 0x5484 */
            {8'h00}, /* 0x5483 */
            {8'h00}, /* 0x5482 */
            {8'h00}, /* 0x5481 */
            {8'h00}, /* 0x5480 */
            {8'h00}, /* 0x547f */
            {8'h00}, /* 0x547e */
            {8'h00}, /* 0x547d */
            {8'h00}, /* 0x547c */
            {8'h00}, /* 0x547b */
            {8'h00}, /* 0x547a */
            {8'h00}, /* 0x5479 */
            {8'h00}, /* 0x5478 */
            {8'h00}, /* 0x5477 */
            {8'h00}, /* 0x5476 */
            {8'h00}, /* 0x5475 */
            {8'h00}, /* 0x5474 */
            {8'h00}, /* 0x5473 */
            {8'h00}, /* 0x5472 */
            {8'h00}, /* 0x5471 */
            {8'h00}, /* 0x5470 */
            {8'h00}, /* 0x546f */
            {8'h00}, /* 0x546e */
            {8'h00}, /* 0x546d */
            {8'h00}, /* 0x546c */
            {8'h00}, /* 0x546b */
            {8'h00}, /* 0x546a */
            {8'h00}, /* 0x5469 */
            {8'h00}, /* 0x5468 */
            {8'h00}, /* 0x5467 */
            {8'h00}, /* 0x5466 */
            {8'h00}, /* 0x5465 */
            {8'h00}, /* 0x5464 */
            {8'h00}, /* 0x5463 */
            {8'h00}, /* 0x5462 */
            {8'h00}, /* 0x5461 */
            {8'h00}, /* 0x5460 */
            {8'h00}, /* 0x545f */
            {8'h00}, /* 0x545e */
            {8'h00}, /* 0x545d */
            {8'h00}, /* 0x545c */
            {8'h00}, /* 0x545b */
            {8'h00}, /* 0x545a */
            {8'h00}, /* 0x5459 */
            {8'h00}, /* 0x5458 */
            {8'h00}, /* 0x5457 */
            {8'h00}, /* 0x5456 */
            {8'h00}, /* 0x5455 */
            {8'h00}, /* 0x5454 */
            {8'h00}, /* 0x5453 */
            {8'h00}, /* 0x5452 */
            {8'h00}, /* 0x5451 */
            {8'h00}, /* 0x5450 */
            {8'h00}, /* 0x544f */
            {8'h00}, /* 0x544e */
            {8'h00}, /* 0x544d */
            {8'h00}, /* 0x544c */
            {8'h00}, /* 0x544b */
            {8'h00}, /* 0x544a */
            {8'h00}, /* 0x5449 */
            {8'h00}, /* 0x5448 */
            {8'h00}, /* 0x5447 */
            {8'h00}, /* 0x5446 */
            {8'h00}, /* 0x5445 */
            {8'h00}, /* 0x5444 */
            {8'h00}, /* 0x5443 */
            {8'h00}, /* 0x5442 */
            {8'h00}, /* 0x5441 */
            {8'h00}, /* 0x5440 */
            {8'h00}, /* 0x543f */
            {8'h00}, /* 0x543e */
            {8'h00}, /* 0x543d */
            {8'h00}, /* 0x543c */
            {8'h00}, /* 0x543b */
            {8'h00}, /* 0x543a */
            {8'h00}, /* 0x5439 */
            {8'h00}, /* 0x5438 */
            {8'h00}, /* 0x5437 */
            {8'h00}, /* 0x5436 */
            {8'h00}, /* 0x5435 */
            {8'h00}, /* 0x5434 */
            {8'h00}, /* 0x5433 */
            {8'h00}, /* 0x5432 */
            {8'h00}, /* 0x5431 */
            {8'h00}, /* 0x5430 */
            {8'h00}, /* 0x542f */
            {8'h00}, /* 0x542e */
            {8'h00}, /* 0x542d */
            {8'h00}, /* 0x542c */
            {8'h00}, /* 0x542b */
            {8'h00}, /* 0x542a */
            {8'h00}, /* 0x5429 */
            {8'h00}, /* 0x5428 */
            {8'h00}, /* 0x5427 */
            {8'h00}, /* 0x5426 */
            {8'h00}, /* 0x5425 */
            {8'h00}, /* 0x5424 */
            {8'h00}, /* 0x5423 */
            {8'h00}, /* 0x5422 */
            {8'h00}, /* 0x5421 */
            {8'h00}, /* 0x5420 */
            {8'h00}, /* 0x541f */
            {8'h00}, /* 0x541e */
            {8'h00}, /* 0x541d */
            {8'h00}, /* 0x541c */
            {8'h00}, /* 0x541b */
            {8'h00}, /* 0x541a */
            {8'h00}, /* 0x5419 */
            {8'h00}, /* 0x5418 */
            {8'h00}, /* 0x5417 */
            {8'h00}, /* 0x5416 */
            {8'h00}, /* 0x5415 */
            {8'h00}, /* 0x5414 */
            {8'h00}, /* 0x5413 */
            {8'h00}, /* 0x5412 */
            {8'h00}, /* 0x5411 */
            {8'h00}, /* 0x5410 */
            {8'h00}, /* 0x540f */
            {8'h00}, /* 0x540e */
            {8'h00}, /* 0x540d */
            {8'h00}, /* 0x540c */
            {8'h00}, /* 0x540b */
            {8'h00}, /* 0x540a */
            {8'h00}, /* 0x5409 */
            {8'h00}, /* 0x5408 */
            {8'h00}, /* 0x5407 */
            {8'h00}, /* 0x5406 */
            {8'h00}, /* 0x5405 */
            {8'h00}, /* 0x5404 */
            {8'h00}, /* 0x5403 */
            {8'h00}, /* 0x5402 */
            {8'h00}, /* 0x5401 */
            {8'h00}, /* 0x5400 */
            {8'h00}, /* 0x53ff */
            {8'h00}, /* 0x53fe */
            {8'h00}, /* 0x53fd */
            {8'h00}, /* 0x53fc */
            {8'h00}, /* 0x53fb */
            {8'h00}, /* 0x53fa */
            {8'h00}, /* 0x53f9 */
            {8'h00}, /* 0x53f8 */
            {8'h00}, /* 0x53f7 */
            {8'h00}, /* 0x53f6 */
            {8'h00}, /* 0x53f5 */
            {8'h00}, /* 0x53f4 */
            {8'h00}, /* 0x53f3 */
            {8'h00}, /* 0x53f2 */
            {8'h00}, /* 0x53f1 */
            {8'h00}, /* 0x53f0 */
            {8'h00}, /* 0x53ef */
            {8'h00}, /* 0x53ee */
            {8'h00}, /* 0x53ed */
            {8'h00}, /* 0x53ec */
            {8'h00}, /* 0x53eb */
            {8'h00}, /* 0x53ea */
            {8'h00}, /* 0x53e9 */
            {8'h00}, /* 0x53e8 */
            {8'h00}, /* 0x53e7 */
            {8'h00}, /* 0x53e6 */
            {8'h00}, /* 0x53e5 */
            {8'h00}, /* 0x53e4 */
            {8'h00}, /* 0x53e3 */
            {8'h00}, /* 0x53e2 */
            {8'h00}, /* 0x53e1 */
            {8'h00}, /* 0x53e0 */
            {8'h00}, /* 0x53df */
            {8'h00}, /* 0x53de */
            {8'h00}, /* 0x53dd */
            {8'h00}, /* 0x53dc */
            {8'h00}, /* 0x53db */
            {8'h00}, /* 0x53da */
            {8'h00}, /* 0x53d9 */
            {8'h00}, /* 0x53d8 */
            {8'h00}, /* 0x53d7 */
            {8'h00}, /* 0x53d6 */
            {8'h00}, /* 0x53d5 */
            {8'h00}, /* 0x53d4 */
            {8'h00}, /* 0x53d3 */
            {8'h00}, /* 0x53d2 */
            {8'h00}, /* 0x53d1 */
            {8'h00}, /* 0x53d0 */
            {8'h00}, /* 0x53cf */
            {8'h00}, /* 0x53ce */
            {8'h00}, /* 0x53cd */
            {8'h00}, /* 0x53cc */
            {8'h00}, /* 0x53cb */
            {8'h00}, /* 0x53ca */
            {8'h00}, /* 0x53c9 */
            {8'h00}, /* 0x53c8 */
            {8'h00}, /* 0x53c7 */
            {8'h00}, /* 0x53c6 */
            {8'h00}, /* 0x53c5 */
            {8'h00}, /* 0x53c4 */
            {8'h00}, /* 0x53c3 */
            {8'h00}, /* 0x53c2 */
            {8'h00}, /* 0x53c1 */
            {8'h00}, /* 0x53c0 */
            {8'h00}, /* 0x53bf */
            {8'h00}, /* 0x53be */
            {8'h00}, /* 0x53bd */
            {8'h00}, /* 0x53bc */
            {8'h00}, /* 0x53bb */
            {8'h00}, /* 0x53ba */
            {8'h00}, /* 0x53b9 */
            {8'h00}, /* 0x53b8 */
            {8'h00}, /* 0x53b7 */
            {8'h00}, /* 0x53b6 */
            {8'h00}, /* 0x53b5 */
            {8'h00}, /* 0x53b4 */
            {8'h00}, /* 0x53b3 */
            {8'h00}, /* 0x53b2 */
            {8'h00}, /* 0x53b1 */
            {8'h00}, /* 0x53b0 */
            {8'h00}, /* 0x53af */
            {8'h00}, /* 0x53ae */
            {8'h00}, /* 0x53ad */
            {8'h00}, /* 0x53ac */
            {8'h00}, /* 0x53ab */
            {8'h00}, /* 0x53aa */
            {8'h00}, /* 0x53a9 */
            {8'h00}, /* 0x53a8 */
            {8'h00}, /* 0x53a7 */
            {8'h00}, /* 0x53a6 */
            {8'h00}, /* 0x53a5 */
            {8'h00}, /* 0x53a4 */
            {8'h00}, /* 0x53a3 */
            {8'h00}, /* 0x53a2 */
            {8'h00}, /* 0x53a1 */
            {8'h00}, /* 0x53a0 */
            {8'h00}, /* 0x539f */
            {8'h00}, /* 0x539e */
            {8'h00}, /* 0x539d */
            {8'h00}, /* 0x539c */
            {8'h00}, /* 0x539b */
            {8'h00}, /* 0x539a */
            {8'h00}, /* 0x5399 */
            {8'h00}, /* 0x5398 */
            {8'h00}, /* 0x5397 */
            {8'h00}, /* 0x5396 */
            {8'h00}, /* 0x5395 */
            {8'h00}, /* 0x5394 */
            {8'h00}, /* 0x5393 */
            {8'h00}, /* 0x5392 */
            {8'h00}, /* 0x5391 */
            {8'h00}, /* 0x5390 */
            {8'h00}, /* 0x538f */
            {8'h00}, /* 0x538e */
            {8'h00}, /* 0x538d */
            {8'h00}, /* 0x538c */
            {8'h00}, /* 0x538b */
            {8'h00}, /* 0x538a */
            {8'h00}, /* 0x5389 */
            {8'h00}, /* 0x5388 */
            {8'h00}, /* 0x5387 */
            {8'h00}, /* 0x5386 */
            {8'h00}, /* 0x5385 */
            {8'h00}, /* 0x5384 */
            {8'h00}, /* 0x5383 */
            {8'h00}, /* 0x5382 */
            {8'h00}, /* 0x5381 */
            {8'h00}, /* 0x5380 */
            {8'h00}, /* 0x537f */
            {8'h00}, /* 0x537e */
            {8'h00}, /* 0x537d */
            {8'h00}, /* 0x537c */
            {8'h00}, /* 0x537b */
            {8'h00}, /* 0x537a */
            {8'h00}, /* 0x5379 */
            {8'h00}, /* 0x5378 */
            {8'h00}, /* 0x5377 */
            {8'h00}, /* 0x5376 */
            {8'h00}, /* 0x5375 */
            {8'h00}, /* 0x5374 */
            {8'h00}, /* 0x5373 */
            {8'h00}, /* 0x5372 */
            {8'h00}, /* 0x5371 */
            {8'h00}, /* 0x5370 */
            {8'h00}, /* 0x536f */
            {8'h00}, /* 0x536e */
            {8'h00}, /* 0x536d */
            {8'h00}, /* 0x536c */
            {8'h00}, /* 0x536b */
            {8'h00}, /* 0x536a */
            {8'h00}, /* 0x5369 */
            {8'h00}, /* 0x5368 */
            {8'h00}, /* 0x5367 */
            {8'h00}, /* 0x5366 */
            {8'h00}, /* 0x5365 */
            {8'h00}, /* 0x5364 */
            {8'h00}, /* 0x5363 */
            {8'h00}, /* 0x5362 */
            {8'h00}, /* 0x5361 */
            {8'h00}, /* 0x5360 */
            {8'h00}, /* 0x535f */
            {8'h00}, /* 0x535e */
            {8'h00}, /* 0x535d */
            {8'h00}, /* 0x535c */
            {8'h00}, /* 0x535b */
            {8'h00}, /* 0x535a */
            {8'h00}, /* 0x5359 */
            {8'h00}, /* 0x5358 */
            {8'h00}, /* 0x5357 */
            {8'h00}, /* 0x5356 */
            {8'h00}, /* 0x5355 */
            {8'h00}, /* 0x5354 */
            {8'h00}, /* 0x5353 */
            {8'h00}, /* 0x5352 */
            {8'h00}, /* 0x5351 */
            {8'h00}, /* 0x5350 */
            {8'h00}, /* 0x534f */
            {8'h00}, /* 0x534e */
            {8'h00}, /* 0x534d */
            {8'h00}, /* 0x534c */
            {8'h00}, /* 0x534b */
            {8'h00}, /* 0x534a */
            {8'h00}, /* 0x5349 */
            {8'h00}, /* 0x5348 */
            {8'h00}, /* 0x5347 */
            {8'h00}, /* 0x5346 */
            {8'h00}, /* 0x5345 */
            {8'h00}, /* 0x5344 */
            {8'h00}, /* 0x5343 */
            {8'h00}, /* 0x5342 */
            {8'h00}, /* 0x5341 */
            {8'h00}, /* 0x5340 */
            {8'h00}, /* 0x533f */
            {8'h00}, /* 0x533e */
            {8'h00}, /* 0x533d */
            {8'h00}, /* 0x533c */
            {8'h00}, /* 0x533b */
            {8'h00}, /* 0x533a */
            {8'h00}, /* 0x5339 */
            {8'h00}, /* 0x5338 */
            {8'h00}, /* 0x5337 */
            {8'h00}, /* 0x5336 */
            {8'h00}, /* 0x5335 */
            {8'h00}, /* 0x5334 */
            {8'h00}, /* 0x5333 */
            {8'h00}, /* 0x5332 */
            {8'h00}, /* 0x5331 */
            {8'h00}, /* 0x5330 */
            {8'h00}, /* 0x532f */
            {8'h00}, /* 0x532e */
            {8'h00}, /* 0x532d */
            {8'h00}, /* 0x532c */
            {8'h00}, /* 0x532b */
            {8'h00}, /* 0x532a */
            {8'h00}, /* 0x5329 */
            {8'h00}, /* 0x5328 */
            {8'h00}, /* 0x5327 */
            {8'h00}, /* 0x5326 */
            {8'h00}, /* 0x5325 */
            {8'h00}, /* 0x5324 */
            {8'h00}, /* 0x5323 */
            {8'h00}, /* 0x5322 */
            {8'h00}, /* 0x5321 */
            {8'h00}, /* 0x5320 */
            {8'h00}, /* 0x531f */
            {8'h00}, /* 0x531e */
            {8'h00}, /* 0x531d */
            {8'h00}, /* 0x531c */
            {8'h00}, /* 0x531b */
            {8'h00}, /* 0x531a */
            {8'h00}, /* 0x5319 */
            {8'h00}, /* 0x5318 */
            {8'h00}, /* 0x5317 */
            {8'h00}, /* 0x5316 */
            {8'h00}, /* 0x5315 */
            {8'h00}, /* 0x5314 */
            {8'h00}, /* 0x5313 */
            {8'h00}, /* 0x5312 */
            {8'h00}, /* 0x5311 */
            {8'h00}, /* 0x5310 */
            {8'h00}, /* 0x530f */
            {8'h00}, /* 0x530e */
            {8'h00}, /* 0x530d */
            {8'h00}, /* 0x530c */
            {8'h00}, /* 0x530b */
            {8'h00}, /* 0x530a */
            {8'h00}, /* 0x5309 */
            {8'h00}, /* 0x5308 */
            {8'h00}, /* 0x5307 */
            {8'h00}, /* 0x5306 */
            {8'h00}, /* 0x5305 */
            {8'h00}, /* 0x5304 */
            {8'h00}, /* 0x5303 */
            {8'h00}, /* 0x5302 */
            {8'h00}, /* 0x5301 */
            {8'h00}, /* 0x5300 */
            {8'h00}, /* 0x52ff */
            {8'h00}, /* 0x52fe */
            {8'h00}, /* 0x52fd */
            {8'h00}, /* 0x52fc */
            {8'h00}, /* 0x52fb */
            {8'h00}, /* 0x52fa */
            {8'h00}, /* 0x52f9 */
            {8'h00}, /* 0x52f8 */
            {8'h00}, /* 0x52f7 */
            {8'h00}, /* 0x52f6 */
            {8'h00}, /* 0x52f5 */
            {8'h00}, /* 0x52f4 */
            {8'h00}, /* 0x52f3 */
            {8'h00}, /* 0x52f2 */
            {8'h00}, /* 0x52f1 */
            {8'h00}, /* 0x52f0 */
            {8'h00}, /* 0x52ef */
            {8'h00}, /* 0x52ee */
            {8'h00}, /* 0x52ed */
            {8'h00}, /* 0x52ec */
            {8'h00}, /* 0x52eb */
            {8'h00}, /* 0x52ea */
            {8'h00}, /* 0x52e9 */
            {8'h00}, /* 0x52e8 */
            {8'h00}, /* 0x52e7 */
            {8'h00}, /* 0x52e6 */
            {8'h00}, /* 0x52e5 */
            {8'h00}, /* 0x52e4 */
            {8'h00}, /* 0x52e3 */
            {8'h00}, /* 0x52e2 */
            {8'h00}, /* 0x52e1 */
            {8'h00}, /* 0x52e0 */
            {8'h00}, /* 0x52df */
            {8'h00}, /* 0x52de */
            {8'h00}, /* 0x52dd */
            {8'h00}, /* 0x52dc */
            {8'h00}, /* 0x52db */
            {8'h00}, /* 0x52da */
            {8'h00}, /* 0x52d9 */
            {8'h00}, /* 0x52d8 */
            {8'h00}, /* 0x52d7 */
            {8'h00}, /* 0x52d6 */
            {8'h00}, /* 0x52d5 */
            {8'h00}, /* 0x52d4 */
            {8'h00}, /* 0x52d3 */
            {8'h00}, /* 0x52d2 */
            {8'h00}, /* 0x52d1 */
            {8'h00}, /* 0x52d0 */
            {8'h00}, /* 0x52cf */
            {8'h00}, /* 0x52ce */
            {8'h00}, /* 0x52cd */
            {8'h00}, /* 0x52cc */
            {8'h00}, /* 0x52cb */
            {8'h00}, /* 0x52ca */
            {8'h00}, /* 0x52c9 */
            {8'h00}, /* 0x52c8 */
            {8'h00}, /* 0x52c7 */
            {8'h00}, /* 0x52c6 */
            {8'h00}, /* 0x52c5 */
            {8'h00}, /* 0x52c4 */
            {8'h00}, /* 0x52c3 */
            {8'h00}, /* 0x52c2 */
            {8'h00}, /* 0x52c1 */
            {8'h00}, /* 0x52c0 */
            {8'h00}, /* 0x52bf */
            {8'h00}, /* 0x52be */
            {8'h00}, /* 0x52bd */
            {8'h00}, /* 0x52bc */
            {8'h00}, /* 0x52bb */
            {8'h00}, /* 0x52ba */
            {8'h00}, /* 0x52b9 */
            {8'h00}, /* 0x52b8 */
            {8'h00}, /* 0x52b7 */
            {8'h00}, /* 0x52b6 */
            {8'h00}, /* 0x52b5 */
            {8'h00}, /* 0x52b4 */
            {8'h00}, /* 0x52b3 */
            {8'h00}, /* 0x52b2 */
            {8'h00}, /* 0x52b1 */
            {8'h00}, /* 0x52b0 */
            {8'h00}, /* 0x52af */
            {8'h00}, /* 0x52ae */
            {8'h00}, /* 0x52ad */
            {8'h00}, /* 0x52ac */
            {8'h00}, /* 0x52ab */
            {8'h00}, /* 0x52aa */
            {8'h00}, /* 0x52a9 */
            {8'h00}, /* 0x52a8 */
            {8'h00}, /* 0x52a7 */
            {8'h00}, /* 0x52a6 */
            {8'h00}, /* 0x52a5 */
            {8'h00}, /* 0x52a4 */
            {8'h00}, /* 0x52a3 */
            {8'h00}, /* 0x52a2 */
            {8'h00}, /* 0x52a1 */
            {8'h00}, /* 0x52a0 */
            {8'h00}, /* 0x529f */
            {8'h00}, /* 0x529e */
            {8'h00}, /* 0x529d */
            {8'h00}, /* 0x529c */
            {8'h00}, /* 0x529b */
            {8'h00}, /* 0x529a */
            {8'h00}, /* 0x5299 */
            {8'h00}, /* 0x5298 */
            {8'h00}, /* 0x5297 */
            {8'h00}, /* 0x5296 */
            {8'h00}, /* 0x5295 */
            {8'h00}, /* 0x5294 */
            {8'h00}, /* 0x5293 */
            {8'h00}, /* 0x5292 */
            {8'h00}, /* 0x5291 */
            {8'h00}, /* 0x5290 */
            {8'h00}, /* 0x528f */
            {8'h00}, /* 0x528e */
            {8'h00}, /* 0x528d */
            {8'h00}, /* 0x528c */
            {8'h00}, /* 0x528b */
            {8'h00}, /* 0x528a */
            {8'h00}, /* 0x5289 */
            {8'h00}, /* 0x5288 */
            {8'h00}, /* 0x5287 */
            {8'h00}, /* 0x5286 */
            {8'h00}, /* 0x5285 */
            {8'h00}, /* 0x5284 */
            {8'h00}, /* 0x5283 */
            {8'h00}, /* 0x5282 */
            {8'h00}, /* 0x5281 */
            {8'h00}, /* 0x5280 */
            {8'h00}, /* 0x527f */
            {8'h00}, /* 0x527e */
            {8'h00}, /* 0x527d */
            {8'h00}, /* 0x527c */
            {8'h00}, /* 0x527b */
            {8'h00}, /* 0x527a */
            {8'h00}, /* 0x5279 */
            {8'h00}, /* 0x5278 */
            {8'h00}, /* 0x5277 */
            {8'h00}, /* 0x5276 */
            {8'h00}, /* 0x5275 */
            {8'h00}, /* 0x5274 */
            {8'h00}, /* 0x5273 */
            {8'h00}, /* 0x5272 */
            {8'h00}, /* 0x5271 */
            {8'h00}, /* 0x5270 */
            {8'h00}, /* 0x526f */
            {8'h00}, /* 0x526e */
            {8'h00}, /* 0x526d */
            {8'h00}, /* 0x526c */
            {8'h00}, /* 0x526b */
            {8'h00}, /* 0x526a */
            {8'h00}, /* 0x5269 */
            {8'h00}, /* 0x5268 */
            {8'h00}, /* 0x5267 */
            {8'h00}, /* 0x5266 */
            {8'h00}, /* 0x5265 */
            {8'h00}, /* 0x5264 */
            {8'h00}, /* 0x5263 */
            {8'h00}, /* 0x5262 */
            {8'h00}, /* 0x5261 */
            {8'h00}, /* 0x5260 */
            {8'h00}, /* 0x525f */
            {8'h00}, /* 0x525e */
            {8'h00}, /* 0x525d */
            {8'h00}, /* 0x525c */
            {8'h00}, /* 0x525b */
            {8'h00}, /* 0x525a */
            {8'h00}, /* 0x5259 */
            {8'h00}, /* 0x5258 */
            {8'h00}, /* 0x5257 */
            {8'h00}, /* 0x5256 */
            {8'h00}, /* 0x5255 */
            {8'h00}, /* 0x5254 */
            {8'h00}, /* 0x5253 */
            {8'h00}, /* 0x5252 */
            {8'h00}, /* 0x5251 */
            {8'h00}, /* 0x5250 */
            {8'h00}, /* 0x524f */
            {8'h00}, /* 0x524e */
            {8'h00}, /* 0x524d */
            {8'h00}, /* 0x524c */
            {8'h00}, /* 0x524b */
            {8'h00}, /* 0x524a */
            {8'h00}, /* 0x5249 */
            {8'h00}, /* 0x5248 */
            {8'h00}, /* 0x5247 */
            {8'h00}, /* 0x5246 */
            {8'h00}, /* 0x5245 */
            {8'h00}, /* 0x5244 */
            {8'h00}, /* 0x5243 */
            {8'h00}, /* 0x5242 */
            {8'h00}, /* 0x5241 */
            {8'h00}, /* 0x5240 */
            {8'h00}, /* 0x523f */
            {8'h00}, /* 0x523e */
            {8'h00}, /* 0x523d */
            {8'h00}, /* 0x523c */
            {8'h00}, /* 0x523b */
            {8'h00}, /* 0x523a */
            {8'h00}, /* 0x5239 */
            {8'h00}, /* 0x5238 */
            {8'h00}, /* 0x5237 */
            {8'h00}, /* 0x5236 */
            {8'h00}, /* 0x5235 */
            {8'h00}, /* 0x5234 */
            {8'h00}, /* 0x5233 */
            {8'h00}, /* 0x5232 */
            {8'h00}, /* 0x5231 */
            {8'h00}, /* 0x5230 */
            {8'h00}, /* 0x522f */
            {8'h00}, /* 0x522e */
            {8'h00}, /* 0x522d */
            {8'h00}, /* 0x522c */
            {8'h00}, /* 0x522b */
            {8'h00}, /* 0x522a */
            {8'h00}, /* 0x5229 */
            {8'h00}, /* 0x5228 */
            {8'h00}, /* 0x5227 */
            {8'h00}, /* 0x5226 */
            {8'h00}, /* 0x5225 */
            {8'h00}, /* 0x5224 */
            {8'h00}, /* 0x5223 */
            {8'h00}, /* 0x5222 */
            {8'h00}, /* 0x5221 */
            {8'h00}, /* 0x5220 */
            {8'h00}, /* 0x521f */
            {8'h00}, /* 0x521e */
            {8'h00}, /* 0x521d */
            {8'h00}, /* 0x521c */
            {8'h00}, /* 0x521b */
            {8'h00}, /* 0x521a */
            {8'h00}, /* 0x5219 */
            {8'h00}, /* 0x5218 */
            {8'h00}, /* 0x5217 */
            {8'h00}, /* 0x5216 */
            {8'h00}, /* 0x5215 */
            {8'h00}, /* 0x5214 */
            {8'h00}, /* 0x5213 */
            {8'h00}, /* 0x5212 */
            {8'h00}, /* 0x5211 */
            {8'h00}, /* 0x5210 */
            {8'h00}, /* 0x520f */
            {8'h00}, /* 0x520e */
            {8'h00}, /* 0x520d */
            {8'h00}, /* 0x520c */
            {8'h00}, /* 0x520b */
            {8'h00}, /* 0x520a */
            {8'h00}, /* 0x5209 */
            {8'h00}, /* 0x5208 */
            {8'h00}, /* 0x5207 */
            {8'h00}, /* 0x5206 */
            {8'h00}, /* 0x5205 */
            {8'h00}, /* 0x5204 */
            {8'h00}, /* 0x5203 */
            {8'h00}, /* 0x5202 */
            {8'h00}, /* 0x5201 */
            {8'h00}, /* 0x5200 */
            {8'h00}, /* 0x51ff */
            {8'h00}, /* 0x51fe */
            {8'h00}, /* 0x51fd */
            {8'h00}, /* 0x51fc */
            {8'h00}, /* 0x51fb */
            {8'h00}, /* 0x51fa */
            {8'h00}, /* 0x51f9 */
            {8'h00}, /* 0x51f8 */
            {8'h00}, /* 0x51f7 */
            {8'h00}, /* 0x51f6 */
            {8'h00}, /* 0x51f5 */
            {8'h00}, /* 0x51f4 */
            {8'h00}, /* 0x51f3 */
            {8'h00}, /* 0x51f2 */
            {8'h00}, /* 0x51f1 */
            {8'h00}, /* 0x51f0 */
            {8'h00}, /* 0x51ef */
            {8'h00}, /* 0x51ee */
            {8'h00}, /* 0x51ed */
            {8'h00}, /* 0x51ec */
            {8'h00}, /* 0x51eb */
            {8'h00}, /* 0x51ea */
            {8'h00}, /* 0x51e9 */
            {8'h00}, /* 0x51e8 */
            {8'h00}, /* 0x51e7 */
            {8'h00}, /* 0x51e6 */
            {8'h00}, /* 0x51e5 */
            {8'h00}, /* 0x51e4 */
            {8'h00}, /* 0x51e3 */
            {8'h00}, /* 0x51e2 */
            {8'h00}, /* 0x51e1 */
            {8'h00}, /* 0x51e0 */
            {8'h00}, /* 0x51df */
            {8'h00}, /* 0x51de */
            {8'h00}, /* 0x51dd */
            {8'h00}, /* 0x51dc */
            {8'h00}, /* 0x51db */
            {8'h00}, /* 0x51da */
            {8'h00}, /* 0x51d9 */
            {8'h00}, /* 0x51d8 */
            {8'h00}, /* 0x51d7 */
            {8'h00}, /* 0x51d6 */
            {8'h00}, /* 0x51d5 */
            {8'h00}, /* 0x51d4 */
            {8'h00}, /* 0x51d3 */
            {8'h00}, /* 0x51d2 */
            {8'h00}, /* 0x51d1 */
            {8'h00}, /* 0x51d0 */
            {8'h00}, /* 0x51cf */
            {8'h00}, /* 0x51ce */
            {8'h00}, /* 0x51cd */
            {8'h00}, /* 0x51cc */
            {8'h00}, /* 0x51cb */
            {8'h00}, /* 0x51ca */
            {8'h00}, /* 0x51c9 */
            {8'h00}, /* 0x51c8 */
            {8'h00}, /* 0x51c7 */
            {8'h00}, /* 0x51c6 */
            {8'h00}, /* 0x51c5 */
            {8'h00}, /* 0x51c4 */
            {8'h00}, /* 0x51c3 */
            {8'h00}, /* 0x51c2 */
            {8'h00}, /* 0x51c1 */
            {8'h00}, /* 0x51c0 */
            {8'h00}, /* 0x51bf */
            {8'h00}, /* 0x51be */
            {8'h00}, /* 0x51bd */
            {8'h00}, /* 0x51bc */
            {8'h00}, /* 0x51bb */
            {8'h00}, /* 0x51ba */
            {8'h00}, /* 0x51b9 */
            {8'h00}, /* 0x51b8 */
            {8'h00}, /* 0x51b7 */
            {8'h00}, /* 0x51b6 */
            {8'h00}, /* 0x51b5 */
            {8'h00}, /* 0x51b4 */
            {8'h00}, /* 0x51b3 */
            {8'h00}, /* 0x51b2 */
            {8'h00}, /* 0x51b1 */
            {8'h00}, /* 0x51b0 */
            {8'h00}, /* 0x51af */
            {8'h00}, /* 0x51ae */
            {8'h00}, /* 0x51ad */
            {8'h00}, /* 0x51ac */
            {8'h00}, /* 0x51ab */
            {8'h00}, /* 0x51aa */
            {8'h00}, /* 0x51a9 */
            {8'h00}, /* 0x51a8 */
            {8'h00}, /* 0x51a7 */
            {8'h00}, /* 0x51a6 */
            {8'h00}, /* 0x51a5 */
            {8'h00}, /* 0x51a4 */
            {8'h00}, /* 0x51a3 */
            {8'h00}, /* 0x51a2 */
            {8'h00}, /* 0x51a1 */
            {8'h00}, /* 0x51a0 */
            {8'h00}, /* 0x519f */
            {8'h00}, /* 0x519e */
            {8'h00}, /* 0x519d */
            {8'h00}, /* 0x519c */
            {8'h00}, /* 0x519b */
            {8'h00}, /* 0x519a */
            {8'h00}, /* 0x5199 */
            {8'h00}, /* 0x5198 */
            {8'h00}, /* 0x5197 */
            {8'h00}, /* 0x5196 */
            {8'h00}, /* 0x5195 */
            {8'h00}, /* 0x5194 */
            {8'h00}, /* 0x5193 */
            {8'h00}, /* 0x5192 */
            {8'h00}, /* 0x5191 */
            {8'h00}, /* 0x5190 */
            {8'h00}, /* 0x518f */
            {8'h00}, /* 0x518e */
            {8'h00}, /* 0x518d */
            {8'h00}, /* 0x518c */
            {8'h00}, /* 0x518b */
            {8'h00}, /* 0x518a */
            {8'h00}, /* 0x5189 */
            {8'h00}, /* 0x5188 */
            {8'h00}, /* 0x5187 */
            {8'h00}, /* 0x5186 */
            {8'h00}, /* 0x5185 */
            {8'h00}, /* 0x5184 */
            {8'h00}, /* 0x5183 */
            {8'h00}, /* 0x5182 */
            {8'h00}, /* 0x5181 */
            {8'h00}, /* 0x5180 */
            {8'h00}, /* 0x517f */
            {8'h00}, /* 0x517e */
            {8'h00}, /* 0x517d */
            {8'h00}, /* 0x517c */
            {8'h00}, /* 0x517b */
            {8'h00}, /* 0x517a */
            {8'h00}, /* 0x5179 */
            {8'h00}, /* 0x5178 */
            {8'h00}, /* 0x5177 */
            {8'h00}, /* 0x5176 */
            {8'h00}, /* 0x5175 */
            {8'h00}, /* 0x5174 */
            {8'h00}, /* 0x5173 */
            {8'h00}, /* 0x5172 */
            {8'h00}, /* 0x5171 */
            {8'h00}, /* 0x5170 */
            {8'h00}, /* 0x516f */
            {8'h00}, /* 0x516e */
            {8'h00}, /* 0x516d */
            {8'h00}, /* 0x516c */
            {8'h00}, /* 0x516b */
            {8'h00}, /* 0x516a */
            {8'h00}, /* 0x5169 */
            {8'h00}, /* 0x5168 */
            {8'h00}, /* 0x5167 */
            {8'h00}, /* 0x5166 */
            {8'h00}, /* 0x5165 */
            {8'h00}, /* 0x5164 */
            {8'h00}, /* 0x5163 */
            {8'h00}, /* 0x5162 */
            {8'h00}, /* 0x5161 */
            {8'h00}, /* 0x5160 */
            {8'h00}, /* 0x515f */
            {8'h00}, /* 0x515e */
            {8'h00}, /* 0x515d */
            {8'h00}, /* 0x515c */
            {8'h00}, /* 0x515b */
            {8'h00}, /* 0x515a */
            {8'h00}, /* 0x5159 */
            {8'h00}, /* 0x5158 */
            {8'h00}, /* 0x5157 */
            {8'h00}, /* 0x5156 */
            {8'h00}, /* 0x5155 */
            {8'h00}, /* 0x5154 */
            {8'h00}, /* 0x5153 */
            {8'h00}, /* 0x5152 */
            {8'h00}, /* 0x5151 */
            {8'h00}, /* 0x5150 */
            {8'h00}, /* 0x514f */
            {8'h00}, /* 0x514e */
            {8'h00}, /* 0x514d */
            {8'h00}, /* 0x514c */
            {8'h00}, /* 0x514b */
            {8'h00}, /* 0x514a */
            {8'h00}, /* 0x5149 */
            {8'h00}, /* 0x5148 */
            {8'h00}, /* 0x5147 */
            {8'h00}, /* 0x5146 */
            {8'h00}, /* 0x5145 */
            {8'h00}, /* 0x5144 */
            {8'h00}, /* 0x5143 */
            {8'h00}, /* 0x5142 */
            {8'h00}, /* 0x5141 */
            {8'h00}, /* 0x5140 */
            {8'h00}, /* 0x513f */
            {8'h00}, /* 0x513e */
            {8'h00}, /* 0x513d */
            {8'h00}, /* 0x513c */
            {8'h00}, /* 0x513b */
            {8'h00}, /* 0x513a */
            {8'h00}, /* 0x5139 */
            {8'h00}, /* 0x5138 */
            {8'h00}, /* 0x5137 */
            {8'h00}, /* 0x5136 */
            {8'h00}, /* 0x5135 */
            {8'h00}, /* 0x5134 */
            {8'h00}, /* 0x5133 */
            {8'h00}, /* 0x5132 */
            {8'h00}, /* 0x5131 */
            {8'h00}, /* 0x5130 */
            {8'h00}, /* 0x512f */
            {8'h00}, /* 0x512e */
            {8'h00}, /* 0x512d */
            {8'h00}, /* 0x512c */
            {8'h00}, /* 0x512b */
            {8'h00}, /* 0x512a */
            {8'h00}, /* 0x5129 */
            {8'h00}, /* 0x5128 */
            {8'h00}, /* 0x5127 */
            {8'h00}, /* 0x5126 */
            {8'h00}, /* 0x5125 */
            {8'h00}, /* 0x5124 */
            {8'h00}, /* 0x5123 */
            {8'h00}, /* 0x5122 */
            {8'h00}, /* 0x5121 */
            {8'h00}, /* 0x5120 */
            {8'h00}, /* 0x511f */
            {8'h00}, /* 0x511e */
            {8'h00}, /* 0x511d */
            {8'h00}, /* 0x511c */
            {8'h00}, /* 0x511b */
            {8'h00}, /* 0x511a */
            {8'h00}, /* 0x5119 */
            {8'h00}, /* 0x5118 */
            {8'h00}, /* 0x5117 */
            {8'h00}, /* 0x5116 */
            {8'h00}, /* 0x5115 */
            {8'h00}, /* 0x5114 */
            {8'h00}, /* 0x5113 */
            {8'h00}, /* 0x5112 */
            {8'h00}, /* 0x5111 */
            {8'h00}, /* 0x5110 */
            {8'h00}, /* 0x510f */
            {8'h00}, /* 0x510e */
            {8'h00}, /* 0x510d */
            {8'h00}, /* 0x510c */
            {8'h00}, /* 0x510b */
            {8'h00}, /* 0x510a */
            {8'h00}, /* 0x5109 */
            {8'h00}, /* 0x5108 */
            {8'h00}, /* 0x5107 */
            {8'h00}, /* 0x5106 */
            {8'h00}, /* 0x5105 */
            {8'h00}, /* 0x5104 */
            {8'h00}, /* 0x5103 */
            {8'h00}, /* 0x5102 */
            {8'h00}, /* 0x5101 */
            {8'h00}, /* 0x5100 */
            {8'h00}, /* 0x50ff */
            {8'h00}, /* 0x50fe */
            {8'h00}, /* 0x50fd */
            {8'h00}, /* 0x50fc */
            {8'h00}, /* 0x50fb */
            {8'h00}, /* 0x50fa */
            {8'h00}, /* 0x50f9 */
            {8'h00}, /* 0x50f8 */
            {8'h00}, /* 0x50f7 */
            {8'h00}, /* 0x50f6 */
            {8'h00}, /* 0x50f5 */
            {8'h00}, /* 0x50f4 */
            {8'h00}, /* 0x50f3 */
            {8'h00}, /* 0x50f2 */
            {8'h00}, /* 0x50f1 */
            {8'h00}, /* 0x50f0 */
            {8'h00}, /* 0x50ef */
            {8'h00}, /* 0x50ee */
            {8'h00}, /* 0x50ed */
            {8'h00}, /* 0x50ec */
            {8'h00}, /* 0x50eb */
            {8'h00}, /* 0x50ea */
            {8'h00}, /* 0x50e9 */
            {8'h00}, /* 0x50e8 */
            {8'h00}, /* 0x50e7 */
            {8'h00}, /* 0x50e6 */
            {8'h00}, /* 0x50e5 */
            {8'h00}, /* 0x50e4 */
            {8'h00}, /* 0x50e3 */
            {8'h00}, /* 0x50e2 */
            {8'h00}, /* 0x50e1 */
            {8'h00}, /* 0x50e0 */
            {8'h00}, /* 0x50df */
            {8'h00}, /* 0x50de */
            {8'h00}, /* 0x50dd */
            {8'h00}, /* 0x50dc */
            {8'h00}, /* 0x50db */
            {8'h00}, /* 0x50da */
            {8'h00}, /* 0x50d9 */
            {8'h00}, /* 0x50d8 */
            {8'h00}, /* 0x50d7 */
            {8'h00}, /* 0x50d6 */
            {8'h00}, /* 0x50d5 */
            {8'h00}, /* 0x50d4 */
            {8'h00}, /* 0x50d3 */
            {8'h00}, /* 0x50d2 */
            {8'h00}, /* 0x50d1 */
            {8'h00}, /* 0x50d0 */
            {8'h00}, /* 0x50cf */
            {8'h00}, /* 0x50ce */
            {8'h00}, /* 0x50cd */
            {8'h00}, /* 0x50cc */
            {8'h00}, /* 0x50cb */
            {8'h00}, /* 0x50ca */
            {8'h00}, /* 0x50c9 */
            {8'h00}, /* 0x50c8 */
            {8'h00}, /* 0x50c7 */
            {8'h00}, /* 0x50c6 */
            {8'h00}, /* 0x50c5 */
            {8'h00}, /* 0x50c4 */
            {8'h00}, /* 0x50c3 */
            {8'h00}, /* 0x50c2 */
            {8'h00}, /* 0x50c1 */
            {8'h00}, /* 0x50c0 */
            {8'h00}, /* 0x50bf */
            {8'h00}, /* 0x50be */
            {8'h00}, /* 0x50bd */
            {8'h00}, /* 0x50bc */
            {8'h00}, /* 0x50bb */
            {8'h00}, /* 0x50ba */
            {8'h00}, /* 0x50b9 */
            {8'h00}, /* 0x50b8 */
            {8'h00}, /* 0x50b7 */
            {8'h00}, /* 0x50b6 */
            {8'h00}, /* 0x50b5 */
            {8'h00}, /* 0x50b4 */
            {8'h00}, /* 0x50b3 */
            {8'h00}, /* 0x50b2 */
            {8'h00}, /* 0x50b1 */
            {8'h00}, /* 0x50b0 */
            {8'h00}, /* 0x50af */
            {8'h00}, /* 0x50ae */
            {8'h00}, /* 0x50ad */
            {8'h00}, /* 0x50ac */
            {8'h00}, /* 0x50ab */
            {8'h00}, /* 0x50aa */
            {8'h00}, /* 0x50a9 */
            {8'h00}, /* 0x50a8 */
            {8'h00}, /* 0x50a7 */
            {8'h00}, /* 0x50a6 */
            {8'h00}, /* 0x50a5 */
            {8'h00}, /* 0x50a4 */
            {8'h00}, /* 0x50a3 */
            {8'h00}, /* 0x50a2 */
            {8'h00}, /* 0x50a1 */
            {8'h00}, /* 0x50a0 */
            {8'h00}, /* 0x509f */
            {8'h00}, /* 0x509e */
            {8'h00}, /* 0x509d */
            {8'h00}, /* 0x509c */
            {8'h00}, /* 0x509b */
            {8'h00}, /* 0x509a */
            {8'h00}, /* 0x5099 */
            {8'h00}, /* 0x5098 */
            {8'h00}, /* 0x5097 */
            {8'h00}, /* 0x5096 */
            {8'h00}, /* 0x5095 */
            {8'h00}, /* 0x5094 */
            {8'h00}, /* 0x5093 */
            {8'h00}, /* 0x5092 */
            {8'h00}, /* 0x5091 */
            {8'h00}, /* 0x5090 */
            {8'h00}, /* 0x508f */
            {8'h00}, /* 0x508e */
            {8'h00}, /* 0x508d */
            {8'h00}, /* 0x508c */
            {8'h00}, /* 0x508b */
            {8'h00}, /* 0x508a */
            {8'h00}, /* 0x5089 */
            {8'h00}, /* 0x5088 */
            {8'h00}, /* 0x5087 */
            {8'h00}, /* 0x5086 */
            {8'h00}, /* 0x5085 */
            {8'h00}, /* 0x5084 */
            {8'h00}, /* 0x5083 */
            {8'h00}, /* 0x5082 */
            {8'h00}, /* 0x5081 */
            {8'h00}, /* 0x5080 */
            {8'h00}, /* 0x507f */
            {8'h00}, /* 0x507e */
            {8'h00}, /* 0x507d */
            {8'h00}, /* 0x507c */
            {8'h00}, /* 0x507b */
            {8'h00}, /* 0x507a */
            {8'h00}, /* 0x5079 */
            {8'h00}, /* 0x5078 */
            {8'h00}, /* 0x5077 */
            {8'h00}, /* 0x5076 */
            {8'h00}, /* 0x5075 */
            {8'h00}, /* 0x5074 */
            {8'h00}, /* 0x5073 */
            {8'h00}, /* 0x5072 */
            {8'h00}, /* 0x5071 */
            {8'h00}, /* 0x5070 */
            {8'h00}, /* 0x506f */
            {8'h00}, /* 0x506e */
            {8'h00}, /* 0x506d */
            {8'h00}, /* 0x506c */
            {8'h00}, /* 0x506b */
            {8'h00}, /* 0x506a */
            {8'h00}, /* 0x5069 */
            {8'h00}, /* 0x5068 */
            {8'h00}, /* 0x5067 */
            {8'h00}, /* 0x5066 */
            {8'h00}, /* 0x5065 */
            {8'h00}, /* 0x5064 */
            {8'h00}, /* 0x5063 */
            {8'h00}, /* 0x5062 */
            {8'h00}, /* 0x5061 */
            {8'h00}, /* 0x5060 */
            {8'h00}, /* 0x505f */
            {8'h00}, /* 0x505e */
            {8'h00}, /* 0x505d */
            {8'h00}, /* 0x505c */
            {8'h00}, /* 0x505b */
            {8'h00}, /* 0x505a */
            {8'h00}, /* 0x5059 */
            {8'h00}, /* 0x5058 */
            {8'h00}, /* 0x5057 */
            {8'h00}, /* 0x5056 */
            {8'h00}, /* 0x5055 */
            {8'h00}, /* 0x5054 */
            {8'h00}, /* 0x5053 */
            {8'h00}, /* 0x5052 */
            {8'h00}, /* 0x5051 */
            {8'h00}, /* 0x5050 */
            {8'h00}, /* 0x504f */
            {8'h00}, /* 0x504e */
            {8'h00}, /* 0x504d */
            {8'h00}, /* 0x504c */
            {8'h00}, /* 0x504b */
            {8'h00}, /* 0x504a */
            {8'h00}, /* 0x5049 */
            {8'h00}, /* 0x5048 */
            {8'h00}, /* 0x5047 */
            {8'h00}, /* 0x5046 */
            {8'h00}, /* 0x5045 */
            {8'h00}, /* 0x5044 */
            {8'h00}, /* 0x5043 */
            {8'h00}, /* 0x5042 */
            {8'h00}, /* 0x5041 */
            {8'h00}, /* 0x5040 */
            {8'h00}, /* 0x503f */
            {8'h00}, /* 0x503e */
            {8'h00}, /* 0x503d */
            {8'h00}, /* 0x503c */
            {8'h00}, /* 0x503b */
            {8'h00}, /* 0x503a */
            {8'h00}, /* 0x5039 */
            {8'h00}, /* 0x5038 */
            {8'h00}, /* 0x5037 */
            {8'h00}, /* 0x5036 */
            {8'h00}, /* 0x5035 */
            {8'h00}, /* 0x5034 */
            {8'h00}, /* 0x5033 */
            {8'h00}, /* 0x5032 */
            {8'h00}, /* 0x5031 */
            {8'h00}, /* 0x5030 */
            {8'h00}, /* 0x502f */
            {8'h00}, /* 0x502e */
            {8'h00}, /* 0x502d */
            {8'h00}, /* 0x502c */
            {8'h00}, /* 0x502b */
            {8'h00}, /* 0x502a */
            {8'h00}, /* 0x5029 */
            {8'h00}, /* 0x5028 */
            {8'h00}, /* 0x5027 */
            {8'h00}, /* 0x5026 */
            {8'h00}, /* 0x5025 */
            {8'h00}, /* 0x5024 */
            {8'h00}, /* 0x5023 */
            {8'h00}, /* 0x5022 */
            {8'h00}, /* 0x5021 */
            {8'h00}, /* 0x5020 */
            {8'h00}, /* 0x501f */
            {8'h00}, /* 0x501e */
            {8'h00}, /* 0x501d */
            {8'h00}, /* 0x501c */
            {8'h00}, /* 0x501b */
            {8'h00}, /* 0x501a */
            {8'h00}, /* 0x5019 */
            {8'h00}, /* 0x5018 */
            {8'h00}, /* 0x5017 */
            {8'h00}, /* 0x5016 */
            {8'h00}, /* 0x5015 */
            {8'h00}, /* 0x5014 */
            {8'h00}, /* 0x5013 */
            {8'h00}, /* 0x5012 */
            {8'h00}, /* 0x5011 */
            {8'h00}, /* 0x5010 */
            {8'h00}, /* 0x500f */
            {8'h00}, /* 0x500e */
            {8'h00}, /* 0x500d */
            {8'h00}, /* 0x500c */
            {8'h00}, /* 0x500b */
            {8'h00}, /* 0x500a */
            {8'h00}, /* 0x5009 */
            {8'h00}, /* 0x5008 */
            {8'h00}, /* 0x5007 */
            {8'h00}, /* 0x5006 */
            {8'h00}, /* 0x5005 */
            {8'h00}, /* 0x5004 */
            {8'h00}, /* 0x5003 */
            {8'h00}, /* 0x5002 */
            {8'h00}, /* 0x5001 */
            {8'h00}, /* 0x5000 */
            {8'h00}, /* 0x4fff */
            {8'h00}, /* 0x4ffe */
            {8'h00}, /* 0x4ffd */
            {8'h00}, /* 0x4ffc */
            {8'h00}, /* 0x4ffb */
            {8'h00}, /* 0x4ffa */
            {8'h00}, /* 0x4ff9 */
            {8'h00}, /* 0x4ff8 */
            {8'h00}, /* 0x4ff7 */
            {8'h00}, /* 0x4ff6 */
            {8'h00}, /* 0x4ff5 */
            {8'h00}, /* 0x4ff4 */
            {8'h00}, /* 0x4ff3 */
            {8'h00}, /* 0x4ff2 */
            {8'h00}, /* 0x4ff1 */
            {8'h00}, /* 0x4ff0 */
            {8'h00}, /* 0x4fef */
            {8'h00}, /* 0x4fee */
            {8'h00}, /* 0x4fed */
            {8'h00}, /* 0x4fec */
            {8'h00}, /* 0x4feb */
            {8'h00}, /* 0x4fea */
            {8'h00}, /* 0x4fe9 */
            {8'h00}, /* 0x4fe8 */
            {8'h00}, /* 0x4fe7 */
            {8'h00}, /* 0x4fe6 */
            {8'h00}, /* 0x4fe5 */
            {8'h00}, /* 0x4fe4 */
            {8'h00}, /* 0x4fe3 */
            {8'h00}, /* 0x4fe2 */
            {8'h00}, /* 0x4fe1 */
            {8'h00}, /* 0x4fe0 */
            {8'h00}, /* 0x4fdf */
            {8'h00}, /* 0x4fde */
            {8'h00}, /* 0x4fdd */
            {8'h00}, /* 0x4fdc */
            {8'h00}, /* 0x4fdb */
            {8'h00}, /* 0x4fda */
            {8'h00}, /* 0x4fd9 */
            {8'h00}, /* 0x4fd8 */
            {8'h00}, /* 0x4fd7 */
            {8'h00}, /* 0x4fd6 */
            {8'h00}, /* 0x4fd5 */
            {8'h00}, /* 0x4fd4 */
            {8'h00}, /* 0x4fd3 */
            {8'h00}, /* 0x4fd2 */
            {8'h00}, /* 0x4fd1 */
            {8'h00}, /* 0x4fd0 */
            {8'h00}, /* 0x4fcf */
            {8'h00}, /* 0x4fce */
            {8'h00}, /* 0x4fcd */
            {8'h00}, /* 0x4fcc */
            {8'h00}, /* 0x4fcb */
            {8'h00}, /* 0x4fca */
            {8'h00}, /* 0x4fc9 */
            {8'h00}, /* 0x4fc8 */
            {8'h00}, /* 0x4fc7 */
            {8'h00}, /* 0x4fc6 */
            {8'h00}, /* 0x4fc5 */
            {8'h00}, /* 0x4fc4 */
            {8'h00}, /* 0x4fc3 */
            {8'h00}, /* 0x4fc2 */
            {8'h00}, /* 0x4fc1 */
            {8'h00}, /* 0x4fc0 */
            {8'h00}, /* 0x4fbf */
            {8'h00}, /* 0x4fbe */
            {8'h00}, /* 0x4fbd */
            {8'h00}, /* 0x4fbc */
            {8'h00}, /* 0x4fbb */
            {8'h00}, /* 0x4fba */
            {8'h00}, /* 0x4fb9 */
            {8'h00}, /* 0x4fb8 */
            {8'h00}, /* 0x4fb7 */
            {8'h00}, /* 0x4fb6 */
            {8'h00}, /* 0x4fb5 */
            {8'h00}, /* 0x4fb4 */
            {8'h00}, /* 0x4fb3 */
            {8'h00}, /* 0x4fb2 */
            {8'h00}, /* 0x4fb1 */
            {8'h00}, /* 0x4fb0 */
            {8'h00}, /* 0x4faf */
            {8'h00}, /* 0x4fae */
            {8'h00}, /* 0x4fad */
            {8'h00}, /* 0x4fac */
            {8'h00}, /* 0x4fab */
            {8'h00}, /* 0x4faa */
            {8'h00}, /* 0x4fa9 */
            {8'h00}, /* 0x4fa8 */
            {8'h00}, /* 0x4fa7 */
            {8'h00}, /* 0x4fa6 */
            {8'h00}, /* 0x4fa5 */
            {8'h00}, /* 0x4fa4 */
            {8'h00}, /* 0x4fa3 */
            {8'h00}, /* 0x4fa2 */
            {8'h00}, /* 0x4fa1 */
            {8'h00}, /* 0x4fa0 */
            {8'h00}, /* 0x4f9f */
            {8'h00}, /* 0x4f9e */
            {8'h00}, /* 0x4f9d */
            {8'h00}, /* 0x4f9c */
            {8'h00}, /* 0x4f9b */
            {8'h00}, /* 0x4f9a */
            {8'h00}, /* 0x4f99 */
            {8'h00}, /* 0x4f98 */
            {8'h00}, /* 0x4f97 */
            {8'h00}, /* 0x4f96 */
            {8'h00}, /* 0x4f95 */
            {8'h00}, /* 0x4f94 */
            {8'h00}, /* 0x4f93 */
            {8'h00}, /* 0x4f92 */
            {8'h00}, /* 0x4f91 */
            {8'h00}, /* 0x4f90 */
            {8'h00}, /* 0x4f8f */
            {8'h00}, /* 0x4f8e */
            {8'h00}, /* 0x4f8d */
            {8'h00}, /* 0x4f8c */
            {8'h00}, /* 0x4f8b */
            {8'h00}, /* 0x4f8a */
            {8'h00}, /* 0x4f89 */
            {8'h00}, /* 0x4f88 */
            {8'h00}, /* 0x4f87 */
            {8'h00}, /* 0x4f86 */
            {8'h00}, /* 0x4f85 */
            {8'h00}, /* 0x4f84 */
            {8'h00}, /* 0x4f83 */
            {8'h00}, /* 0x4f82 */
            {8'h00}, /* 0x4f81 */
            {8'h00}, /* 0x4f80 */
            {8'h00}, /* 0x4f7f */
            {8'h00}, /* 0x4f7e */
            {8'h00}, /* 0x4f7d */
            {8'h00}, /* 0x4f7c */
            {8'h00}, /* 0x4f7b */
            {8'h00}, /* 0x4f7a */
            {8'h00}, /* 0x4f79 */
            {8'h00}, /* 0x4f78 */
            {8'h00}, /* 0x4f77 */
            {8'h00}, /* 0x4f76 */
            {8'h00}, /* 0x4f75 */
            {8'h00}, /* 0x4f74 */
            {8'h00}, /* 0x4f73 */
            {8'h00}, /* 0x4f72 */
            {8'h00}, /* 0x4f71 */
            {8'h00}, /* 0x4f70 */
            {8'h00}, /* 0x4f6f */
            {8'h00}, /* 0x4f6e */
            {8'h00}, /* 0x4f6d */
            {8'h00}, /* 0x4f6c */
            {8'h00}, /* 0x4f6b */
            {8'h00}, /* 0x4f6a */
            {8'h00}, /* 0x4f69 */
            {8'h00}, /* 0x4f68 */
            {8'h00}, /* 0x4f67 */
            {8'h00}, /* 0x4f66 */
            {8'h00}, /* 0x4f65 */
            {8'h00}, /* 0x4f64 */
            {8'h00}, /* 0x4f63 */
            {8'h00}, /* 0x4f62 */
            {8'h00}, /* 0x4f61 */
            {8'h00}, /* 0x4f60 */
            {8'h00}, /* 0x4f5f */
            {8'h00}, /* 0x4f5e */
            {8'h00}, /* 0x4f5d */
            {8'h00}, /* 0x4f5c */
            {8'h00}, /* 0x4f5b */
            {8'h00}, /* 0x4f5a */
            {8'h00}, /* 0x4f59 */
            {8'h00}, /* 0x4f58 */
            {8'h00}, /* 0x4f57 */
            {8'h00}, /* 0x4f56 */
            {8'h00}, /* 0x4f55 */
            {8'h00}, /* 0x4f54 */
            {8'h00}, /* 0x4f53 */
            {8'h00}, /* 0x4f52 */
            {8'h00}, /* 0x4f51 */
            {8'h00}, /* 0x4f50 */
            {8'h00}, /* 0x4f4f */
            {8'h00}, /* 0x4f4e */
            {8'h00}, /* 0x4f4d */
            {8'h00}, /* 0x4f4c */
            {8'h00}, /* 0x4f4b */
            {8'h00}, /* 0x4f4a */
            {8'h00}, /* 0x4f49 */
            {8'h00}, /* 0x4f48 */
            {8'h00}, /* 0x4f47 */
            {8'h00}, /* 0x4f46 */
            {8'h00}, /* 0x4f45 */
            {8'h00}, /* 0x4f44 */
            {8'h00}, /* 0x4f43 */
            {8'h00}, /* 0x4f42 */
            {8'h00}, /* 0x4f41 */
            {8'h00}, /* 0x4f40 */
            {8'h00}, /* 0x4f3f */
            {8'h00}, /* 0x4f3e */
            {8'h00}, /* 0x4f3d */
            {8'h00}, /* 0x4f3c */
            {8'h00}, /* 0x4f3b */
            {8'h00}, /* 0x4f3a */
            {8'h00}, /* 0x4f39 */
            {8'h00}, /* 0x4f38 */
            {8'h00}, /* 0x4f37 */
            {8'h00}, /* 0x4f36 */
            {8'h00}, /* 0x4f35 */
            {8'h00}, /* 0x4f34 */
            {8'h00}, /* 0x4f33 */
            {8'h00}, /* 0x4f32 */
            {8'h00}, /* 0x4f31 */
            {8'h00}, /* 0x4f30 */
            {8'h00}, /* 0x4f2f */
            {8'h00}, /* 0x4f2e */
            {8'h00}, /* 0x4f2d */
            {8'h00}, /* 0x4f2c */
            {8'h00}, /* 0x4f2b */
            {8'h00}, /* 0x4f2a */
            {8'h00}, /* 0x4f29 */
            {8'h00}, /* 0x4f28 */
            {8'h00}, /* 0x4f27 */
            {8'h00}, /* 0x4f26 */
            {8'h00}, /* 0x4f25 */
            {8'h00}, /* 0x4f24 */
            {8'h00}, /* 0x4f23 */
            {8'h00}, /* 0x4f22 */
            {8'h00}, /* 0x4f21 */
            {8'h00}, /* 0x4f20 */
            {8'h00}, /* 0x4f1f */
            {8'h00}, /* 0x4f1e */
            {8'h00}, /* 0x4f1d */
            {8'h00}, /* 0x4f1c */
            {8'h00}, /* 0x4f1b */
            {8'h00}, /* 0x4f1a */
            {8'h00}, /* 0x4f19 */
            {8'h00}, /* 0x4f18 */
            {8'h00}, /* 0x4f17 */
            {8'h00}, /* 0x4f16 */
            {8'h00}, /* 0x4f15 */
            {8'h00}, /* 0x4f14 */
            {8'h00}, /* 0x4f13 */
            {8'h00}, /* 0x4f12 */
            {8'h00}, /* 0x4f11 */
            {8'h00}, /* 0x4f10 */
            {8'h00}, /* 0x4f0f */
            {8'h00}, /* 0x4f0e */
            {8'h00}, /* 0x4f0d */
            {8'h00}, /* 0x4f0c */
            {8'h00}, /* 0x4f0b */
            {8'h00}, /* 0x4f0a */
            {8'h00}, /* 0x4f09 */
            {8'h00}, /* 0x4f08 */
            {8'h00}, /* 0x4f07 */
            {8'h00}, /* 0x4f06 */
            {8'h00}, /* 0x4f05 */
            {8'h00}, /* 0x4f04 */
            {8'h00}, /* 0x4f03 */
            {8'h00}, /* 0x4f02 */
            {8'h00}, /* 0x4f01 */
            {8'h00}, /* 0x4f00 */
            {8'h00}, /* 0x4eff */
            {8'h00}, /* 0x4efe */
            {8'h00}, /* 0x4efd */
            {8'h00}, /* 0x4efc */
            {8'h00}, /* 0x4efb */
            {8'h00}, /* 0x4efa */
            {8'h00}, /* 0x4ef9 */
            {8'h00}, /* 0x4ef8 */
            {8'h00}, /* 0x4ef7 */
            {8'h00}, /* 0x4ef6 */
            {8'h00}, /* 0x4ef5 */
            {8'h00}, /* 0x4ef4 */
            {8'h00}, /* 0x4ef3 */
            {8'h00}, /* 0x4ef2 */
            {8'h00}, /* 0x4ef1 */
            {8'h00}, /* 0x4ef0 */
            {8'h00}, /* 0x4eef */
            {8'h00}, /* 0x4eee */
            {8'h00}, /* 0x4eed */
            {8'h00}, /* 0x4eec */
            {8'h00}, /* 0x4eeb */
            {8'h00}, /* 0x4eea */
            {8'h00}, /* 0x4ee9 */
            {8'h00}, /* 0x4ee8 */
            {8'h00}, /* 0x4ee7 */
            {8'h00}, /* 0x4ee6 */
            {8'h00}, /* 0x4ee5 */
            {8'h00}, /* 0x4ee4 */
            {8'h00}, /* 0x4ee3 */
            {8'h00}, /* 0x4ee2 */
            {8'h00}, /* 0x4ee1 */
            {8'h00}, /* 0x4ee0 */
            {8'h00}, /* 0x4edf */
            {8'h00}, /* 0x4ede */
            {8'h00}, /* 0x4edd */
            {8'h00}, /* 0x4edc */
            {8'h00}, /* 0x4edb */
            {8'h00}, /* 0x4eda */
            {8'h00}, /* 0x4ed9 */
            {8'h00}, /* 0x4ed8 */
            {8'h00}, /* 0x4ed7 */
            {8'h00}, /* 0x4ed6 */
            {8'h00}, /* 0x4ed5 */
            {8'h00}, /* 0x4ed4 */
            {8'h00}, /* 0x4ed3 */
            {8'h00}, /* 0x4ed2 */
            {8'h00}, /* 0x4ed1 */
            {8'h00}, /* 0x4ed0 */
            {8'h00}, /* 0x4ecf */
            {8'h00}, /* 0x4ece */
            {8'h00}, /* 0x4ecd */
            {8'h00}, /* 0x4ecc */
            {8'h00}, /* 0x4ecb */
            {8'h00}, /* 0x4eca */
            {8'h00}, /* 0x4ec9 */
            {8'h00}, /* 0x4ec8 */
            {8'h00}, /* 0x4ec7 */
            {8'h00}, /* 0x4ec6 */
            {8'h00}, /* 0x4ec5 */
            {8'h00}, /* 0x4ec4 */
            {8'h00}, /* 0x4ec3 */
            {8'h00}, /* 0x4ec2 */
            {8'h00}, /* 0x4ec1 */
            {8'h00}, /* 0x4ec0 */
            {8'h00}, /* 0x4ebf */
            {8'h00}, /* 0x4ebe */
            {8'h00}, /* 0x4ebd */
            {8'h00}, /* 0x4ebc */
            {8'h00}, /* 0x4ebb */
            {8'h00}, /* 0x4eba */
            {8'h00}, /* 0x4eb9 */
            {8'h00}, /* 0x4eb8 */
            {8'h00}, /* 0x4eb7 */
            {8'h00}, /* 0x4eb6 */
            {8'h00}, /* 0x4eb5 */
            {8'h00}, /* 0x4eb4 */
            {8'h00}, /* 0x4eb3 */
            {8'h00}, /* 0x4eb2 */
            {8'h00}, /* 0x4eb1 */
            {8'h00}, /* 0x4eb0 */
            {8'h00}, /* 0x4eaf */
            {8'h00}, /* 0x4eae */
            {8'h00}, /* 0x4ead */
            {8'h00}, /* 0x4eac */
            {8'h00}, /* 0x4eab */
            {8'h00}, /* 0x4eaa */
            {8'h00}, /* 0x4ea9 */
            {8'h00}, /* 0x4ea8 */
            {8'h00}, /* 0x4ea7 */
            {8'h00}, /* 0x4ea6 */
            {8'h00}, /* 0x4ea5 */
            {8'h00}, /* 0x4ea4 */
            {8'h00}, /* 0x4ea3 */
            {8'h00}, /* 0x4ea2 */
            {8'h00}, /* 0x4ea1 */
            {8'h00}, /* 0x4ea0 */
            {8'h00}, /* 0x4e9f */
            {8'h00}, /* 0x4e9e */
            {8'h00}, /* 0x4e9d */
            {8'h00}, /* 0x4e9c */
            {8'h00}, /* 0x4e9b */
            {8'h00}, /* 0x4e9a */
            {8'h00}, /* 0x4e99 */
            {8'h00}, /* 0x4e98 */
            {8'h00}, /* 0x4e97 */
            {8'h00}, /* 0x4e96 */
            {8'h00}, /* 0x4e95 */
            {8'h00}, /* 0x4e94 */
            {8'h00}, /* 0x4e93 */
            {8'h00}, /* 0x4e92 */
            {8'h00}, /* 0x4e91 */
            {8'h00}, /* 0x4e90 */
            {8'h00}, /* 0x4e8f */
            {8'h00}, /* 0x4e8e */
            {8'h00}, /* 0x4e8d */
            {8'h00}, /* 0x4e8c */
            {8'h00}, /* 0x4e8b */
            {8'h00}, /* 0x4e8a */
            {8'h00}, /* 0x4e89 */
            {8'h00}, /* 0x4e88 */
            {8'h00}, /* 0x4e87 */
            {8'h00}, /* 0x4e86 */
            {8'h00}, /* 0x4e85 */
            {8'h00}, /* 0x4e84 */
            {8'h00}, /* 0x4e83 */
            {8'h00}, /* 0x4e82 */
            {8'h00}, /* 0x4e81 */
            {8'h00}, /* 0x4e80 */
            {8'h00}, /* 0x4e7f */
            {8'h00}, /* 0x4e7e */
            {8'h00}, /* 0x4e7d */
            {8'h00}, /* 0x4e7c */
            {8'h00}, /* 0x4e7b */
            {8'h00}, /* 0x4e7a */
            {8'h00}, /* 0x4e79 */
            {8'h00}, /* 0x4e78 */
            {8'h00}, /* 0x4e77 */
            {8'h00}, /* 0x4e76 */
            {8'h00}, /* 0x4e75 */
            {8'h00}, /* 0x4e74 */
            {8'h00}, /* 0x4e73 */
            {8'h00}, /* 0x4e72 */
            {8'h00}, /* 0x4e71 */
            {8'h00}, /* 0x4e70 */
            {8'h00}, /* 0x4e6f */
            {8'h00}, /* 0x4e6e */
            {8'h00}, /* 0x4e6d */
            {8'h00}, /* 0x4e6c */
            {8'h00}, /* 0x4e6b */
            {8'h00}, /* 0x4e6a */
            {8'h00}, /* 0x4e69 */
            {8'h00}, /* 0x4e68 */
            {8'h00}, /* 0x4e67 */
            {8'h00}, /* 0x4e66 */
            {8'h00}, /* 0x4e65 */
            {8'h00}, /* 0x4e64 */
            {8'h00}, /* 0x4e63 */
            {8'h00}, /* 0x4e62 */
            {8'h00}, /* 0x4e61 */
            {8'h00}, /* 0x4e60 */
            {8'h00}, /* 0x4e5f */
            {8'h00}, /* 0x4e5e */
            {8'h00}, /* 0x4e5d */
            {8'h00}, /* 0x4e5c */
            {8'h00}, /* 0x4e5b */
            {8'h00}, /* 0x4e5a */
            {8'h00}, /* 0x4e59 */
            {8'h00}, /* 0x4e58 */
            {8'h00}, /* 0x4e57 */
            {8'h00}, /* 0x4e56 */
            {8'h00}, /* 0x4e55 */
            {8'h00}, /* 0x4e54 */
            {8'h00}, /* 0x4e53 */
            {8'h00}, /* 0x4e52 */
            {8'h00}, /* 0x4e51 */
            {8'h00}, /* 0x4e50 */
            {8'h00}, /* 0x4e4f */
            {8'h00}, /* 0x4e4e */
            {8'h00}, /* 0x4e4d */
            {8'h00}, /* 0x4e4c */
            {8'h00}, /* 0x4e4b */
            {8'h00}, /* 0x4e4a */
            {8'h00}, /* 0x4e49 */
            {8'h00}, /* 0x4e48 */
            {8'h00}, /* 0x4e47 */
            {8'h00}, /* 0x4e46 */
            {8'h00}, /* 0x4e45 */
            {8'h00}, /* 0x4e44 */
            {8'h00}, /* 0x4e43 */
            {8'h00}, /* 0x4e42 */
            {8'h00}, /* 0x4e41 */
            {8'h00}, /* 0x4e40 */
            {8'h00}, /* 0x4e3f */
            {8'h00}, /* 0x4e3e */
            {8'h00}, /* 0x4e3d */
            {8'h00}, /* 0x4e3c */
            {8'h00}, /* 0x4e3b */
            {8'h00}, /* 0x4e3a */
            {8'h00}, /* 0x4e39 */
            {8'h00}, /* 0x4e38 */
            {8'h00}, /* 0x4e37 */
            {8'h00}, /* 0x4e36 */
            {8'h00}, /* 0x4e35 */
            {8'h00}, /* 0x4e34 */
            {8'h00}, /* 0x4e33 */
            {8'h00}, /* 0x4e32 */
            {8'h00}, /* 0x4e31 */
            {8'h00}, /* 0x4e30 */
            {8'h00}, /* 0x4e2f */
            {8'h00}, /* 0x4e2e */
            {8'h00}, /* 0x4e2d */
            {8'h00}, /* 0x4e2c */
            {8'h00}, /* 0x4e2b */
            {8'h00}, /* 0x4e2a */
            {8'h00}, /* 0x4e29 */
            {8'h00}, /* 0x4e28 */
            {8'h00}, /* 0x4e27 */
            {8'h00}, /* 0x4e26 */
            {8'h00}, /* 0x4e25 */
            {8'h00}, /* 0x4e24 */
            {8'h00}, /* 0x4e23 */
            {8'h00}, /* 0x4e22 */
            {8'h00}, /* 0x4e21 */
            {8'h00}, /* 0x4e20 */
            {8'h00}, /* 0x4e1f */
            {8'h00}, /* 0x4e1e */
            {8'h00}, /* 0x4e1d */
            {8'h00}, /* 0x4e1c */
            {8'h00}, /* 0x4e1b */
            {8'h00}, /* 0x4e1a */
            {8'h00}, /* 0x4e19 */
            {8'h00}, /* 0x4e18 */
            {8'h00}, /* 0x4e17 */
            {8'h00}, /* 0x4e16 */
            {8'h00}, /* 0x4e15 */
            {8'h00}, /* 0x4e14 */
            {8'h00}, /* 0x4e13 */
            {8'h00}, /* 0x4e12 */
            {8'h00}, /* 0x4e11 */
            {8'h00}, /* 0x4e10 */
            {8'h00}, /* 0x4e0f */
            {8'h00}, /* 0x4e0e */
            {8'h00}, /* 0x4e0d */
            {8'h00}, /* 0x4e0c */
            {8'h00}, /* 0x4e0b */
            {8'h00}, /* 0x4e0a */
            {8'h00}, /* 0x4e09 */
            {8'h00}, /* 0x4e08 */
            {8'h00}, /* 0x4e07 */
            {8'h00}, /* 0x4e06 */
            {8'h00}, /* 0x4e05 */
            {8'h00}, /* 0x4e04 */
            {8'h00}, /* 0x4e03 */
            {8'h00}, /* 0x4e02 */
            {8'h00}, /* 0x4e01 */
            {8'h00}, /* 0x4e00 */
            {8'h00}, /* 0x4dff */
            {8'h00}, /* 0x4dfe */
            {8'h00}, /* 0x4dfd */
            {8'h00}, /* 0x4dfc */
            {8'h00}, /* 0x4dfb */
            {8'h00}, /* 0x4dfa */
            {8'h00}, /* 0x4df9 */
            {8'h00}, /* 0x4df8 */
            {8'h00}, /* 0x4df7 */
            {8'h00}, /* 0x4df6 */
            {8'h00}, /* 0x4df5 */
            {8'h00}, /* 0x4df4 */
            {8'h00}, /* 0x4df3 */
            {8'h00}, /* 0x4df2 */
            {8'h00}, /* 0x4df1 */
            {8'h00}, /* 0x4df0 */
            {8'h00}, /* 0x4def */
            {8'h00}, /* 0x4dee */
            {8'h00}, /* 0x4ded */
            {8'h00}, /* 0x4dec */
            {8'h00}, /* 0x4deb */
            {8'h00}, /* 0x4dea */
            {8'h00}, /* 0x4de9 */
            {8'h00}, /* 0x4de8 */
            {8'h00}, /* 0x4de7 */
            {8'h00}, /* 0x4de6 */
            {8'h00}, /* 0x4de5 */
            {8'h00}, /* 0x4de4 */
            {8'h00}, /* 0x4de3 */
            {8'h00}, /* 0x4de2 */
            {8'h00}, /* 0x4de1 */
            {8'h00}, /* 0x4de0 */
            {8'h00}, /* 0x4ddf */
            {8'h00}, /* 0x4dde */
            {8'h00}, /* 0x4ddd */
            {8'h00}, /* 0x4ddc */
            {8'h00}, /* 0x4ddb */
            {8'h00}, /* 0x4dda */
            {8'h00}, /* 0x4dd9 */
            {8'h00}, /* 0x4dd8 */
            {8'h00}, /* 0x4dd7 */
            {8'h00}, /* 0x4dd6 */
            {8'h00}, /* 0x4dd5 */
            {8'h00}, /* 0x4dd4 */
            {8'h00}, /* 0x4dd3 */
            {8'h00}, /* 0x4dd2 */
            {8'h00}, /* 0x4dd1 */
            {8'h00}, /* 0x4dd0 */
            {8'h00}, /* 0x4dcf */
            {8'h00}, /* 0x4dce */
            {8'h00}, /* 0x4dcd */
            {8'h00}, /* 0x4dcc */
            {8'h00}, /* 0x4dcb */
            {8'h00}, /* 0x4dca */
            {8'h00}, /* 0x4dc9 */
            {8'h00}, /* 0x4dc8 */
            {8'h00}, /* 0x4dc7 */
            {8'h00}, /* 0x4dc6 */
            {8'h00}, /* 0x4dc5 */
            {8'h00}, /* 0x4dc4 */
            {8'h00}, /* 0x4dc3 */
            {8'h00}, /* 0x4dc2 */
            {8'h00}, /* 0x4dc1 */
            {8'h00}, /* 0x4dc0 */
            {8'h00}, /* 0x4dbf */
            {8'h00}, /* 0x4dbe */
            {8'h00}, /* 0x4dbd */
            {8'h00}, /* 0x4dbc */
            {8'h00}, /* 0x4dbb */
            {8'h00}, /* 0x4dba */
            {8'h00}, /* 0x4db9 */
            {8'h00}, /* 0x4db8 */
            {8'h00}, /* 0x4db7 */
            {8'h00}, /* 0x4db6 */
            {8'h00}, /* 0x4db5 */
            {8'h00}, /* 0x4db4 */
            {8'h00}, /* 0x4db3 */
            {8'h00}, /* 0x4db2 */
            {8'h00}, /* 0x4db1 */
            {8'h00}, /* 0x4db0 */
            {8'h00}, /* 0x4daf */
            {8'h00}, /* 0x4dae */
            {8'h00}, /* 0x4dad */
            {8'h00}, /* 0x4dac */
            {8'h00}, /* 0x4dab */
            {8'h00}, /* 0x4daa */
            {8'h00}, /* 0x4da9 */
            {8'h00}, /* 0x4da8 */
            {8'h00}, /* 0x4da7 */
            {8'h00}, /* 0x4da6 */
            {8'h00}, /* 0x4da5 */
            {8'h00}, /* 0x4da4 */
            {8'h00}, /* 0x4da3 */
            {8'h00}, /* 0x4da2 */
            {8'h00}, /* 0x4da1 */
            {8'h00}, /* 0x4da0 */
            {8'h00}, /* 0x4d9f */
            {8'h00}, /* 0x4d9e */
            {8'h00}, /* 0x4d9d */
            {8'h00}, /* 0x4d9c */
            {8'h00}, /* 0x4d9b */
            {8'h00}, /* 0x4d9a */
            {8'h00}, /* 0x4d99 */
            {8'h00}, /* 0x4d98 */
            {8'h00}, /* 0x4d97 */
            {8'h00}, /* 0x4d96 */
            {8'h00}, /* 0x4d95 */
            {8'h00}, /* 0x4d94 */
            {8'h00}, /* 0x4d93 */
            {8'h00}, /* 0x4d92 */
            {8'h00}, /* 0x4d91 */
            {8'h00}, /* 0x4d90 */
            {8'h00}, /* 0x4d8f */
            {8'h00}, /* 0x4d8e */
            {8'h00}, /* 0x4d8d */
            {8'h00}, /* 0x4d8c */
            {8'h00}, /* 0x4d8b */
            {8'h00}, /* 0x4d8a */
            {8'h00}, /* 0x4d89 */
            {8'h00}, /* 0x4d88 */
            {8'h00}, /* 0x4d87 */
            {8'h00}, /* 0x4d86 */
            {8'h00}, /* 0x4d85 */
            {8'h00}, /* 0x4d84 */
            {8'h00}, /* 0x4d83 */
            {8'h00}, /* 0x4d82 */
            {8'h00}, /* 0x4d81 */
            {8'h00}, /* 0x4d80 */
            {8'h00}, /* 0x4d7f */
            {8'h00}, /* 0x4d7e */
            {8'h00}, /* 0x4d7d */
            {8'h00}, /* 0x4d7c */
            {8'h00}, /* 0x4d7b */
            {8'h00}, /* 0x4d7a */
            {8'h00}, /* 0x4d79 */
            {8'h00}, /* 0x4d78 */
            {8'h00}, /* 0x4d77 */
            {8'h00}, /* 0x4d76 */
            {8'h00}, /* 0x4d75 */
            {8'h00}, /* 0x4d74 */
            {8'h00}, /* 0x4d73 */
            {8'h00}, /* 0x4d72 */
            {8'h00}, /* 0x4d71 */
            {8'h00}, /* 0x4d70 */
            {8'h00}, /* 0x4d6f */
            {8'h00}, /* 0x4d6e */
            {8'h00}, /* 0x4d6d */
            {8'h00}, /* 0x4d6c */
            {8'h00}, /* 0x4d6b */
            {8'h00}, /* 0x4d6a */
            {8'h00}, /* 0x4d69 */
            {8'h00}, /* 0x4d68 */
            {8'h00}, /* 0x4d67 */
            {8'h00}, /* 0x4d66 */
            {8'h00}, /* 0x4d65 */
            {8'h00}, /* 0x4d64 */
            {8'h00}, /* 0x4d63 */
            {8'h00}, /* 0x4d62 */
            {8'h00}, /* 0x4d61 */
            {8'h00}, /* 0x4d60 */
            {8'h00}, /* 0x4d5f */
            {8'h00}, /* 0x4d5e */
            {8'h00}, /* 0x4d5d */
            {8'h00}, /* 0x4d5c */
            {8'h00}, /* 0x4d5b */
            {8'h00}, /* 0x4d5a */
            {8'h00}, /* 0x4d59 */
            {8'h00}, /* 0x4d58 */
            {8'h00}, /* 0x4d57 */
            {8'h00}, /* 0x4d56 */
            {8'h00}, /* 0x4d55 */
            {8'h00}, /* 0x4d54 */
            {8'h00}, /* 0x4d53 */
            {8'h00}, /* 0x4d52 */
            {8'h00}, /* 0x4d51 */
            {8'h00}, /* 0x4d50 */
            {8'h00}, /* 0x4d4f */
            {8'h00}, /* 0x4d4e */
            {8'h00}, /* 0x4d4d */
            {8'h00}, /* 0x4d4c */
            {8'h00}, /* 0x4d4b */
            {8'h00}, /* 0x4d4a */
            {8'h00}, /* 0x4d49 */
            {8'h00}, /* 0x4d48 */
            {8'h00}, /* 0x4d47 */
            {8'h00}, /* 0x4d46 */
            {8'h00}, /* 0x4d45 */
            {8'h00}, /* 0x4d44 */
            {8'h00}, /* 0x4d43 */
            {8'h00}, /* 0x4d42 */
            {8'h00}, /* 0x4d41 */
            {8'h00}, /* 0x4d40 */
            {8'h00}, /* 0x4d3f */
            {8'h00}, /* 0x4d3e */
            {8'h00}, /* 0x4d3d */
            {8'h00}, /* 0x4d3c */
            {8'h00}, /* 0x4d3b */
            {8'h00}, /* 0x4d3a */
            {8'h00}, /* 0x4d39 */
            {8'h00}, /* 0x4d38 */
            {8'h00}, /* 0x4d37 */
            {8'h00}, /* 0x4d36 */
            {8'h00}, /* 0x4d35 */
            {8'h00}, /* 0x4d34 */
            {8'h00}, /* 0x4d33 */
            {8'h00}, /* 0x4d32 */
            {8'h00}, /* 0x4d31 */
            {8'h00}, /* 0x4d30 */
            {8'h00}, /* 0x4d2f */
            {8'h00}, /* 0x4d2e */
            {8'h00}, /* 0x4d2d */
            {8'h00}, /* 0x4d2c */
            {8'h00}, /* 0x4d2b */
            {8'h00}, /* 0x4d2a */
            {8'h00}, /* 0x4d29 */
            {8'h00}, /* 0x4d28 */
            {8'h00}, /* 0x4d27 */
            {8'h00}, /* 0x4d26 */
            {8'h00}, /* 0x4d25 */
            {8'h00}, /* 0x4d24 */
            {8'h00}, /* 0x4d23 */
            {8'h00}, /* 0x4d22 */
            {8'h00}, /* 0x4d21 */
            {8'h00}, /* 0x4d20 */
            {8'h00}, /* 0x4d1f */
            {8'h00}, /* 0x4d1e */
            {8'h00}, /* 0x4d1d */
            {8'h00}, /* 0x4d1c */
            {8'h00}, /* 0x4d1b */
            {8'h00}, /* 0x4d1a */
            {8'h00}, /* 0x4d19 */
            {8'h00}, /* 0x4d18 */
            {8'h00}, /* 0x4d17 */
            {8'h00}, /* 0x4d16 */
            {8'h00}, /* 0x4d15 */
            {8'h00}, /* 0x4d14 */
            {8'h00}, /* 0x4d13 */
            {8'h00}, /* 0x4d12 */
            {8'h00}, /* 0x4d11 */
            {8'h00}, /* 0x4d10 */
            {8'h00}, /* 0x4d0f */
            {8'h00}, /* 0x4d0e */
            {8'h00}, /* 0x4d0d */
            {8'h00}, /* 0x4d0c */
            {8'h00}, /* 0x4d0b */
            {8'h00}, /* 0x4d0a */
            {8'h00}, /* 0x4d09 */
            {8'h00}, /* 0x4d08 */
            {8'h00}, /* 0x4d07 */
            {8'h00}, /* 0x4d06 */
            {8'h00}, /* 0x4d05 */
            {8'h00}, /* 0x4d04 */
            {8'h00}, /* 0x4d03 */
            {8'h00}, /* 0x4d02 */
            {8'h00}, /* 0x4d01 */
            {8'h00}, /* 0x4d00 */
            {8'h00}, /* 0x4cff */
            {8'h00}, /* 0x4cfe */
            {8'h00}, /* 0x4cfd */
            {8'h00}, /* 0x4cfc */
            {8'h00}, /* 0x4cfb */
            {8'h00}, /* 0x4cfa */
            {8'h00}, /* 0x4cf9 */
            {8'h00}, /* 0x4cf8 */
            {8'h00}, /* 0x4cf7 */
            {8'h00}, /* 0x4cf6 */
            {8'h00}, /* 0x4cf5 */
            {8'h00}, /* 0x4cf4 */
            {8'h00}, /* 0x4cf3 */
            {8'h00}, /* 0x4cf2 */
            {8'h00}, /* 0x4cf1 */
            {8'h00}, /* 0x4cf0 */
            {8'h00}, /* 0x4cef */
            {8'h00}, /* 0x4cee */
            {8'h00}, /* 0x4ced */
            {8'h00}, /* 0x4cec */
            {8'h00}, /* 0x4ceb */
            {8'h00}, /* 0x4cea */
            {8'h00}, /* 0x4ce9 */
            {8'h00}, /* 0x4ce8 */
            {8'h00}, /* 0x4ce7 */
            {8'h00}, /* 0x4ce6 */
            {8'h00}, /* 0x4ce5 */
            {8'h00}, /* 0x4ce4 */
            {8'h00}, /* 0x4ce3 */
            {8'h00}, /* 0x4ce2 */
            {8'h00}, /* 0x4ce1 */
            {8'h00}, /* 0x4ce0 */
            {8'h00}, /* 0x4cdf */
            {8'h00}, /* 0x4cde */
            {8'h00}, /* 0x4cdd */
            {8'h00}, /* 0x4cdc */
            {8'h00}, /* 0x4cdb */
            {8'h00}, /* 0x4cda */
            {8'h00}, /* 0x4cd9 */
            {8'h00}, /* 0x4cd8 */
            {8'h00}, /* 0x4cd7 */
            {8'h00}, /* 0x4cd6 */
            {8'h00}, /* 0x4cd5 */
            {8'h00}, /* 0x4cd4 */
            {8'h00}, /* 0x4cd3 */
            {8'h00}, /* 0x4cd2 */
            {8'h00}, /* 0x4cd1 */
            {8'h00}, /* 0x4cd0 */
            {8'h00}, /* 0x4ccf */
            {8'h00}, /* 0x4cce */
            {8'h00}, /* 0x4ccd */
            {8'h00}, /* 0x4ccc */
            {8'h00}, /* 0x4ccb */
            {8'h00}, /* 0x4cca */
            {8'h00}, /* 0x4cc9 */
            {8'h00}, /* 0x4cc8 */
            {8'h00}, /* 0x4cc7 */
            {8'h00}, /* 0x4cc6 */
            {8'h00}, /* 0x4cc5 */
            {8'h00}, /* 0x4cc4 */
            {8'h00}, /* 0x4cc3 */
            {8'h00}, /* 0x4cc2 */
            {8'h00}, /* 0x4cc1 */
            {8'h00}, /* 0x4cc0 */
            {8'h00}, /* 0x4cbf */
            {8'h00}, /* 0x4cbe */
            {8'h00}, /* 0x4cbd */
            {8'h00}, /* 0x4cbc */
            {8'h00}, /* 0x4cbb */
            {8'h00}, /* 0x4cba */
            {8'h00}, /* 0x4cb9 */
            {8'h00}, /* 0x4cb8 */
            {8'h00}, /* 0x4cb7 */
            {8'h00}, /* 0x4cb6 */
            {8'h00}, /* 0x4cb5 */
            {8'h00}, /* 0x4cb4 */
            {8'h00}, /* 0x4cb3 */
            {8'h00}, /* 0x4cb2 */
            {8'h00}, /* 0x4cb1 */
            {8'h00}, /* 0x4cb0 */
            {8'h00}, /* 0x4caf */
            {8'h00}, /* 0x4cae */
            {8'h00}, /* 0x4cad */
            {8'h00}, /* 0x4cac */
            {8'h00}, /* 0x4cab */
            {8'h00}, /* 0x4caa */
            {8'h00}, /* 0x4ca9 */
            {8'h00}, /* 0x4ca8 */
            {8'h00}, /* 0x4ca7 */
            {8'h00}, /* 0x4ca6 */
            {8'h00}, /* 0x4ca5 */
            {8'h00}, /* 0x4ca4 */
            {8'h00}, /* 0x4ca3 */
            {8'h00}, /* 0x4ca2 */
            {8'h00}, /* 0x4ca1 */
            {8'h00}, /* 0x4ca0 */
            {8'h00}, /* 0x4c9f */
            {8'h00}, /* 0x4c9e */
            {8'h00}, /* 0x4c9d */
            {8'h00}, /* 0x4c9c */
            {8'h00}, /* 0x4c9b */
            {8'h00}, /* 0x4c9a */
            {8'h00}, /* 0x4c99 */
            {8'h00}, /* 0x4c98 */
            {8'h00}, /* 0x4c97 */
            {8'h00}, /* 0x4c96 */
            {8'h00}, /* 0x4c95 */
            {8'h00}, /* 0x4c94 */
            {8'h00}, /* 0x4c93 */
            {8'h00}, /* 0x4c92 */
            {8'h00}, /* 0x4c91 */
            {8'h00}, /* 0x4c90 */
            {8'h00}, /* 0x4c8f */
            {8'h00}, /* 0x4c8e */
            {8'h00}, /* 0x4c8d */
            {8'h00}, /* 0x4c8c */
            {8'h00}, /* 0x4c8b */
            {8'h00}, /* 0x4c8a */
            {8'h00}, /* 0x4c89 */
            {8'h00}, /* 0x4c88 */
            {8'h00}, /* 0x4c87 */
            {8'h00}, /* 0x4c86 */
            {8'h00}, /* 0x4c85 */
            {8'h00}, /* 0x4c84 */
            {8'h00}, /* 0x4c83 */
            {8'h00}, /* 0x4c82 */
            {8'h00}, /* 0x4c81 */
            {8'h00}, /* 0x4c80 */
            {8'h00}, /* 0x4c7f */
            {8'h00}, /* 0x4c7e */
            {8'h00}, /* 0x4c7d */
            {8'h00}, /* 0x4c7c */
            {8'h00}, /* 0x4c7b */
            {8'h00}, /* 0x4c7a */
            {8'h00}, /* 0x4c79 */
            {8'h00}, /* 0x4c78 */
            {8'h00}, /* 0x4c77 */
            {8'h00}, /* 0x4c76 */
            {8'h00}, /* 0x4c75 */
            {8'h00}, /* 0x4c74 */
            {8'h00}, /* 0x4c73 */
            {8'h00}, /* 0x4c72 */
            {8'h00}, /* 0x4c71 */
            {8'h00}, /* 0x4c70 */
            {8'h00}, /* 0x4c6f */
            {8'h00}, /* 0x4c6e */
            {8'h00}, /* 0x4c6d */
            {8'h00}, /* 0x4c6c */
            {8'h00}, /* 0x4c6b */
            {8'h00}, /* 0x4c6a */
            {8'h00}, /* 0x4c69 */
            {8'h00}, /* 0x4c68 */
            {8'h00}, /* 0x4c67 */
            {8'h00}, /* 0x4c66 */
            {8'h00}, /* 0x4c65 */
            {8'h00}, /* 0x4c64 */
            {8'h00}, /* 0x4c63 */
            {8'h00}, /* 0x4c62 */
            {8'h00}, /* 0x4c61 */
            {8'h00}, /* 0x4c60 */
            {8'h00}, /* 0x4c5f */
            {8'h00}, /* 0x4c5e */
            {8'h00}, /* 0x4c5d */
            {8'h00}, /* 0x4c5c */
            {8'h00}, /* 0x4c5b */
            {8'h00}, /* 0x4c5a */
            {8'h00}, /* 0x4c59 */
            {8'h00}, /* 0x4c58 */
            {8'h00}, /* 0x4c57 */
            {8'h00}, /* 0x4c56 */
            {8'h00}, /* 0x4c55 */
            {8'h00}, /* 0x4c54 */
            {8'h00}, /* 0x4c53 */
            {8'h00}, /* 0x4c52 */
            {8'h00}, /* 0x4c51 */
            {8'h00}, /* 0x4c50 */
            {8'h00}, /* 0x4c4f */
            {8'h00}, /* 0x4c4e */
            {8'h00}, /* 0x4c4d */
            {8'h00}, /* 0x4c4c */
            {8'h00}, /* 0x4c4b */
            {8'h00}, /* 0x4c4a */
            {8'h00}, /* 0x4c49 */
            {8'h00}, /* 0x4c48 */
            {8'h00}, /* 0x4c47 */
            {8'h00}, /* 0x4c46 */
            {8'h00}, /* 0x4c45 */
            {8'h00}, /* 0x4c44 */
            {8'h00}, /* 0x4c43 */
            {8'h00}, /* 0x4c42 */
            {8'h00}, /* 0x4c41 */
            {8'h00}, /* 0x4c40 */
            {8'h00}, /* 0x4c3f */
            {8'h00}, /* 0x4c3e */
            {8'h00}, /* 0x4c3d */
            {8'h00}, /* 0x4c3c */
            {8'h00}, /* 0x4c3b */
            {8'h00}, /* 0x4c3a */
            {8'h00}, /* 0x4c39 */
            {8'h00}, /* 0x4c38 */
            {8'h00}, /* 0x4c37 */
            {8'h00}, /* 0x4c36 */
            {8'h00}, /* 0x4c35 */
            {8'h00}, /* 0x4c34 */
            {8'h00}, /* 0x4c33 */
            {8'h00}, /* 0x4c32 */
            {8'h00}, /* 0x4c31 */
            {8'h00}, /* 0x4c30 */
            {8'h00}, /* 0x4c2f */
            {8'h00}, /* 0x4c2e */
            {8'h00}, /* 0x4c2d */
            {8'h00}, /* 0x4c2c */
            {8'h00}, /* 0x4c2b */
            {8'h00}, /* 0x4c2a */
            {8'h00}, /* 0x4c29 */
            {8'h00}, /* 0x4c28 */
            {8'h00}, /* 0x4c27 */
            {8'h00}, /* 0x4c26 */
            {8'h00}, /* 0x4c25 */
            {8'h00}, /* 0x4c24 */
            {8'h00}, /* 0x4c23 */
            {8'h00}, /* 0x4c22 */
            {8'h00}, /* 0x4c21 */
            {8'h00}, /* 0x4c20 */
            {8'h00}, /* 0x4c1f */
            {8'h00}, /* 0x4c1e */
            {8'h00}, /* 0x4c1d */
            {8'h00}, /* 0x4c1c */
            {8'h00}, /* 0x4c1b */
            {8'h00}, /* 0x4c1a */
            {8'h00}, /* 0x4c19 */
            {8'h00}, /* 0x4c18 */
            {8'h00}, /* 0x4c17 */
            {8'h00}, /* 0x4c16 */
            {8'h00}, /* 0x4c15 */
            {8'h00}, /* 0x4c14 */
            {8'h00}, /* 0x4c13 */
            {8'h00}, /* 0x4c12 */
            {8'h00}, /* 0x4c11 */
            {8'h00}, /* 0x4c10 */
            {8'h00}, /* 0x4c0f */
            {8'h00}, /* 0x4c0e */
            {8'h00}, /* 0x4c0d */
            {8'h00}, /* 0x4c0c */
            {8'h00}, /* 0x4c0b */
            {8'h00}, /* 0x4c0a */
            {8'h00}, /* 0x4c09 */
            {8'h00}, /* 0x4c08 */
            {8'h00}, /* 0x4c07 */
            {8'h00}, /* 0x4c06 */
            {8'h00}, /* 0x4c05 */
            {8'h00}, /* 0x4c04 */
            {8'h00}, /* 0x4c03 */
            {8'h00}, /* 0x4c02 */
            {8'h00}, /* 0x4c01 */
            {8'h00}, /* 0x4c00 */
            {8'h00}, /* 0x4bff */
            {8'h00}, /* 0x4bfe */
            {8'h00}, /* 0x4bfd */
            {8'h00}, /* 0x4bfc */
            {8'h00}, /* 0x4bfb */
            {8'h00}, /* 0x4bfa */
            {8'h00}, /* 0x4bf9 */
            {8'h00}, /* 0x4bf8 */
            {8'h00}, /* 0x4bf7 */
            {8'h00}, /* 0x4bf6 */
            {8'h00}, /* 0x4bf5 */
            {8'h00}, /* 0x4bf4 */
            {8'h00}, /* 0x4bf3 */
            {8'h00}, /* 0x4bf2 */
            {8'h00}, /* 0x4bf1 */
            {8'h00}, /* 0x4bf0 */
            {8'h00}, /* 0x4bef */
            {8'h00}, /* 0x4bee */
            {8'h00}, /* 0x4bed */
            {8'h00}, /* 0x4bec */
            {8'h00}, /* 0x4beb */
            {8'h00}, /* 0x4bea */
            {8'h00}, /* 0x4be9 */
            {8'h00}, /* 0x4be8 */
            {8'h00}, /* 0x4be7 */
            {8'h00}, /* 0x4be6 */
            {8'h00}, /* 0x4be5 */
            {8'h00}, /* 0x4be4 */
            {8'h00}, /* 0x4be3 */
            {8'h00}, /* 0x4be2 */
            {8'h00}, /* 0x4be1 */
            {8'h00}, /* 0x4be0 */
            {8'h00}, /* 0x4bdf */
            {8'h00}, /* 0x4bde */
            {8'h00}, /* 0x4bdd */
            {8'h00}, /* 0x4bdc */
            {8'h00}, /* 0x4bdb */
            {8'h00}, /* 0x4bda */
            {8'h00}, /* 0x4bd9 */
            {8'h00}, /* 0x4bd8 */
            {8'h00}, /* 0x4bd7 */
            {8'h00}, /* 0x4bd6 */
            {8'h00}, /* 0x4bd5 */
            {8'h00}, /* 0x4bd4 */
            {8'h00}, /* 0x4bd3 */
            {8'h00}, /* 0x4bd2 */
            {8'h00}, /* 0x4bd1 */
            {8'h00}, /* 0x4bd0 */
            {8'h00}, /* 0x4bcf */
            {8'h00}, /* 0x4bce */
            {8'h00}, /* 0x4bcd */
            {8'h00}, /* 0x4bcc */
            {8'h00}, /* 0x4bcb */
            {8'h00}, /* 0x4bca */
            {8'h00}, /* 0x4bc9 */
            {8'h00}, /* 0x4bc8 */
            {8'h00}, /* 0x4bc7 */
            {8'h00}, /* 0x4bc6 */
            {8'h00}, /* 0x4bc5 */
            {8'h00}, /* 0x4bc4 */
            {8'h00}, /* 0x4bc3 */
            {8'h00}, /* 0x4bc2 */
            {8'h00}, /* 0x4bc1 */
            {8'h00}, /* 0x4bc0 */
            {8'h00}, /* 0x4bbf */
            {8'h00}, /* 0x4bbe */
            {8'h00}, /* 0x4bbd */
            {8'h00}, /* 0x4bbc */
            {8'h00}, /* 0x4bbb */
            {8'h00}, /* 0x4bba */
            {8'h00}, /* 0x4bb9 */
            {8'h00}, /* 0x4bb8 */
            {8'h00}, /* 0x4bb7 */
            {8'h00}, /* 0x4bb6 */
            {8'h00}, /* 0x4bb5 */
            {8'h00}, /* 0x4bb4 */
            {8'h00}, /* 0x4bb3 */
            {8'h00}, /* 0x4bb2 */
            {8'h00}, /* 0x4bb1 */
            {8'h00}, /* 0x4bb0 */
            {8'h00}, /* 0x4baf */
            {8'h00}, /* 0x4bae */
            {8'h00}, /* 0x4bad */
            {8'h00}, /* 0x4bac */
            {8'h00}, /* 0x4bab */
            {8'h00}, /* 0x4baa */
            {8'h00}, /* 0x4ba9 */
            {8'h00}, /* 0x4ba8 */
            {8'h00}, /* 0x4ba7 */
            {8'h00}, /* 0x4ba6 */
            {8'h00}, /* 0x4ba5 */
            {8'h00}, /* 0x4ba4 */
            {8'h00}, /* 0x4ba3 */
            {8'h00}, /* 0x4ba2 */
            {8'h00}, /* 0x4ba1 */
            {8'h00}, /* 0x4ba0 */
            {8'h00}, /* 0x4b9f */
            {8'h00}, /* 0x4b9e */
            {8'h00}, /* 0x4b9d */
            {8'h00}, /* 0x4b9c */
            {8'h00}, /* 0x4b9b */
            {8'h00}, /* 0x4b9a */
            {8'h00}, /* 0x4b99 */
            {8'h00}, /* 0x4b98 */
            {8'h00}, /* 0x4b97 */
            {8'h00}, /* 0x4b96 */
            {8'h00}, /* 0x4b95 */
            {8'h00}, /* 0x4b94 */
            {8'h00}, /* 0x4b93 */
            {8'h00}, /* 0x4b92 */
            {8'h00}, /* 0x4b91 */
            {8'h00}, /* 0x4b90 */
            {8'h00}, /* 0x4b8f */
            {8'h00}, /* 0x4b8e */
            {8'h00}, /* 0x4b8d */
            {8'h00}, /* 0x4b8c */
            {8'h00}, /* 0x4b8b */
            {8'h00}, /* 0x4b8a */
            {8'h00}, /* 0x4b89 */
            {8'h00}, /* 0x4b88 */
            {8'h00}, /* 0x4b87 */
            {8'h00}, /* 0x4b86 */
            {8'h00}, /* 0x4b85 */
            {8'h00}, /* 0x4b84 */
            {8'h00}, /* 0x4b83 */
            {8'h00}, /* 0x4b82 */
            {8'h00}, /* 0x4b81 */
            {8'h00}, /* 0x4b80 */
            {8'h00}, /* 0x4b7f */
            {8'h00}, /* 0x4b7e */
            {8'h00}, /* 0x4b7d */
            {8'h00}, /* 0x4b7c */
            {8'h00}, /* 0x4b7b */
            {8'h00}, /* 0x4b7a */
            {8'h00}, /* 0x4b79 */
            {8'h00}, /* 0x4b78 */
            {8'h00}, /* 0x4b77 */
            {8'h00}, /* 0x4b76 */
            {8'h00}, /* 0x4b75 */
            {8'h00}, /* 0x4b74 */
            {8'h00}, /* 0x4b73 */
            {8'h00}, /* 0x4b72 */
            {8'h00}, /* 0x4b71 */
            {8'h00}, /* 0x4b70 */
            {8'h00}, /* 0x4b6f */
            {8'h00}, /* 0x4b6e */
            {8'h00}, /* 0x4b6d */
            {8'h00}, /* 0x4b6c */
            {8'h00}, /* 0x4b6b */
            {8'h00}, /* 0x4b6a */
            {8'h00}, /* 0x4b69 */
            {8'h00}, /* 0x4b68 */
            {8'h00}, /* 0x4b67 */
            {8'h00}, /* 0x4b66 */
            {8'h00}, /* 0x4b65 */
            {8'h00}, /* 0x4b64 */
            {8'h00}, /* 0x4b63 */
            {8'h00}, /* 0x4b62 */
            {8'h00}, /* 0x4b61 */
            {8'h00}, /* 0x4b60 */
            {8'h00}, /* 0x4b5f */
            {8'h00}, /* 0x4b5e */
            {8'h00}, /* 0x4b5d */
            {8'h00}, /* 0x4b5c */
            {8'h00}, /* 0x4b5b */
            {8'h00}, /* 0x4b5a */
            {8'h00}, /* 0x4b59 */
            {8'h00}, /* 0x4b58 */
            {8'h00}, /* 0x4b57 */
            {8'h00}, /* 0x4b56 */
            {8'h00}, /* 0x4b55 */
            {8'h00}, /* 0x4b54 */
            {8'h00}, /* 0x4b53 */
            {8'h00}, /* 0x4b52 */
            {8'h00}, /* 0x4b51 */
            {8'h00}, /* 0x4b50 */
            {8'h00}, /* 0x4b4f */
            {8'h00}, /* 0x4b4e */
            {8'h00}, /* 0x4b4d */
            {8'h00}, /* 0x4b4c */
            {8'h00}, /* 0x4b4b */
            {8'h00}, /* 0x4b4a */
            {8'h00}, /* 0x4b49 */
            {8'h00}, /* 0x4b48 */
            {8'h00}, /* 0x4b47 */
            {8'h00}, /* 0x4b46 */
            {8'h00}, /* 0x4b45 */
            {8'h00}, /* 0x4b44 */
            {8'h00}, /* 0x4b43 */
            {8'h00}, /* 0x4b42 */
            {8'h00}, /* 0x4b41 */
            {8'h00}, /* 0x4b40 */
            {8'h00}, /* 0x4b3f */
            {8'h00}, /* 0x4b3e */
            {8'h00}, /* 0x4b3d */
            {8'h00}, /* 0x4b3c */
            {8'h00}, /* 0x4b3b */
            {8'h00}, /* 0x4b3a */
            {8'h00}, /* 0x4b39 */
            {8'h00}, /* 0x4b38 */
            {8'h00}, /* 0x4b37 */
            {8'h00}, /* 0x4b36 */
            {8'h00}, /* 0x4b35 */
            {8'h00}, /* 0x4b34 */
            {8'h00}, /* 0x4b33 */
            {8'h00}, /* 0x4b32 */
            {8'h00}, /* 0x4b31 */
            {8'h00}, /* 0x4b30 */
            {8'h00}, /* 0x4b2f */
            {8'h00}, /* 0x4b2e */
            {8'h00}, /* 0x4b2d */
            {8'h00}, /* 0x4b2c */
            {8'h00}, /* 0x4b2b */
            {8'h00}, /* 0x4b2a */
            {8'h00}, /* 0x4b29 */
            {8'h00}, /* 0x4b28 */
            {8'h00}, /* 0x4b27 */
            {8'h00}, /* 0x4b26 */
            {8'h00}, /* 0x4b25 */
            {8'h00}, /* 0x4b24 */
            {8'h00}, /* 0x4b23 */
            {8'h00}, /* 0x4b22 */
            {8'h00}, /* 0x4b21 */
            {8'h00}, /* 0x4b20 */
            {8'h00}, /* 0x4b1f */
            {8'h00}, /* 0x4b1e */
            {8'h00}, /* 0x4b1d */
            {8'h00}, /* 0x4b1c */
            {8'h00}, /* 0x4b1b */
            {8'h00}, /* 0x4b1a */
            {8'h00}, /* 0x4b19 */
            {8'h00}, /* 0x4b18 */
            {8'h00}, /* 0x4b17 */
            {8'h00}, /* 0x4b16 */
            {8'h00}, /* 0x4b15 */
            {8'h00}, /* 0x4b14 */
            {8'h00}, /* 0x4b13 */
            {8'h00}, /* 0x4b12 */
            {8'h00}, /* 0x4b11 */
            {8'h00}, /* 0x4b10 */
            {8'h00}, /* 0x4b0f */
            {8'h00}, /* 0x4b0e */
            {8'h00}, /* 0x4b0d */
            {8'h00}, /* 0x4b0c */
            {8'h00}, /* 0x4b0b */
            {8'h00}, /* 0x4b0a */
            {8'h00}, /* 0x4b09 */
            {8'h00}, /* 0x4b08 */
            {8'h00}, /* 0x4b07 */
            {8'h00}, /* 0x4b06 */
            {8'h00}, /* 0x4b05 */
            {8'h00}, /* 0x4b04 */
            {8'h00}, /* 0x4b03 */
            {8'h00}, /* 0x4b02 */
            {8'h00}, /* 0x4b01 */
            {8'h00}, /* 0x4b00 */
            {8'h00}, /* 0x4aff */
            {8'h00}, /* 0x4afe */
            {8'h00}, /* 0x4afd */
            {8'h00}, /* 0x4afc */
            {8'h00}, /* 0x4afb */
            {8'h00}, /* 0x4afa */
            {8'h00}, /* 0x4af9 */
            {8'h00}, /* 0x4af8 */
            {8'h00}, /* 0x4af7 */
            {8'h00}, /* 0x4af6 */
            {8'h00}, /* 0x4af5 */
            {8'h00}, /* 0x4af4 */
            {8'h00}, /* 0x4af3 */
            {8'h00}, /* 0x4af2 */
            {8'h00}, /* 0x4af1 */
            {8'h00}, /* 0x4af0 */
            {8'h00}, /* 0x4aef */
            {8'h00}, /* 0x4aee */
            {8'h00}, /* 0x4aed */
            {8'h00}, /* 0x4aec */
            {8'h00}, /* 0x4aeb */
            {8'h00}, /* 0x4aea */
            {8'h00}, /* 0x4ae9 */
            {8'h00}, /* 0x4ae8 */
            {8'h00}, /* 0x4ae7 */
            {8'h00}, /* 0x4ae6 */
            {8'h00}, /* 0x4ae5 */
            {8'h00}, /* 0x4ae4 */
            {8'h00}, /* 0x4ae3 */
            {8'h00}, /* 0x4ae2 */
            {8'h00}, /* 0x4ae1 */
            {8'h00}, /* 0x4ae0 */
            {8'h00}, /* 0x4adf */
            {8'h00}, /* 0x4ade */
            {8'h00}, /* 0x4add */
            {8'h00}, /* 0x4adc */
            {8'h00}, /* 0x4adb */
            {8'h00}, /* 0x4ada */
            {8'h00}, /* 0x4ad9 */
            {8'h00}, /* 0x4ad8 */
            {8'h00}, /* 0x4ad7 */
            {8'h00}, /* 0x4ad6 */
            {8'h00}, /* 0x4ad5 */
            {8'h00}, /* 0x4ad4 */
            {8'h00}, /* 0x4ad3 */
            {8'h00}, /* 0x4ad2 */
            {8'h00}, /* 0x4ad1 */
            {8'h00}, /* 0x4ad0 */
            {8'h00}, /* 0x4acf */
            {8'h00}, /* 0x4ace */
            {8'h00}, /* 0x4acd */
            {8'h00}, /* 0x4acc */
            {8'h00}, /* 0x4acb */
            {8'h00}, /* 0x4aca */
            {8'h00}, /* 0x4ac9 */
            {8'h00}, /* 0x4ac8 */
            {8'h00}, /* 0x4ac7 */
            {8'h00}, /* 0x4ac6 */
            {8'h00}, /* 0x4ac5 */
            {8'h00}, /* 0x4ac4 */
            {8'h00}, /* 0x4ac3 */
            {8'h00}, /* 0x4ac2 */
            {8'h00}, /* 0x4ac1 */
            {8'h00}, /* 0x4ac0 */
            {8'h00}, /* 0x4abf */
            {8'h00}, /* 0x4abe */
            {8'h00}, /* 0x4abd */
            {8'h00}, /* 0x4abc */
            {8'h00}, /* 0x4abb */
            {8'h00}, /* 0x4aba */
            {8'h00}, /* 0x4ab9 */
            {8'h00}, /* 0x4ab8 */
            {8'h00}, /* 0x4ab7 */
            {8'h00}, /* 0x4ab6 */
            {8'h00}, /* 0x4ab5 */
            {8'h00}, /* 0x4ab4 */
            {8'h00}, /* 0x4ab3 */
            {8'h00}, /* 0x4ab2 */
            {8'h00}, /* 0x4ab1 */
            {8'h00}, /* 0x4ab0 */
            {8'h00}, /* 0x4aaf */
            {8'h00}, /* 0x4aae */
            {8'h00}, /* 0x4aad */
            {8'h00}, /* 0x4aac */
            {8'h00}, /* 0x4aab */
            {8'h00}, /* 0x4aaa */
            {8'h00}, /* 0x4aa9 */
            {8'h00}, /* 0x4aa8 */
            {8'h00}, /* 0x4aa7 */
            {8'h00}, /* 0x4aa6 */
            {8'h00}, /* 0x4aa5 */
            {8'h00}, /* 0x4aa4 */
            {8'h00}, /* 0x4aa3 */
            {8'h00}, /* 0x4aa2 */
            {8'h00}, /* 0x4aa1 */
            {8'h00}, /* 0x4aa0 */
            {8'h00}, /* 0x4a9f */
            {8'h00}, /* 0x4a9e */
            {8'h00}, /* 0x4a9d */
            {8'h00}, /* 0x4a9c */
            {8'h00}, /* 0x4a9b */
            {8'h00}, /* 0x4a9a */
            {8'h00}, /* 0x4a99 */
            {8'h00}, /* 0x4a98 */
            {8'h00}, /* 0x4a97 */
            {8'h00}, /* 0x4a96 */
            {8'h00}, /* 0x4a95 */
            {8'h00}, /* 0x4a94 */
            {8'h00}, /* 0x4a93 */
            {8'h00}, /* 0x4a92 */
            {8'h00}, /* 0x4a91 */
            {8'h00}, /* 0x4a90 */
            {8'h00}, /* 0x4a8f */
            {8'h00}, /* 0x4a8e */
            {8'h00}, /* 0x4a8d */
            {8'h00}, /* 0x4a8c */
            {8'h00}, /* 0x4a8b */
            {8'h00}, /* 0x4a8a */
            {8'h00}, /* 0x4a89 */
            {8'h00}, /* 0x4a88 */
            {8'h00}, /* 0x4a87 */
            {8'h00}, /* 0x4a86 */
            {8'h00}, /* 0x4a85 */
            {8'h00}, /* 0x4a84 */
            {8'h00}, /* 0x4a83 */
            {8'h00}, /* 0x4a82 */
            {8'h00}, /* 0x4a81 */
            {8'h00}, /* 0x4a80 */
            {8'h00}, /* 0x4a7f */
            {8'h00}, /* 0x4a7e */
            {8'h00}, /* 0x4a7d */
            {8'h00}, /* 0x4a7c */
            {8'h00}, /* 0x4a7b */
            {8'h00}, /* 0x4a7a */
            {8'h00}, /* 0x4a79 */
            {8'h00}, /* 0x4a78 */
            {8'h00}, /* 0x4a77 */
            {8'h00}, /* 0x4a76 */
            {8'h00}, /* 0x4a75 */
            {8'h00}, /* 0x4a74 */
            {8'h00}, /* 0x4a73 */
            {8'h00}, /* 0x4a72 */
            {8'h00}, /* 0x4a71 */
            {8'h00}, /* 0x4a70 */
            {8'h00}, /* 0x4a6f */
            {8'h00}, /* 0x4a6e */
            {8'h00}, /* 0x4a6d */
            {8'h00}, /* 0x4a6c */
            {8'h00}, /* 0x4a6b */
            {8'h00}, /* 0x4a6a */
            {8'h00}, /* 0x4a69 */
            {8'h00}, /* 0x4a68 */
            {8'h00}, /* 0x4a67 */
            {8'h00}, /* 0x4a66 */
            {8'h00}, /* 0x4a65 */
            {8'h00}, /* 0x4a64 */
            {8'h00}, /* 0x4a63 */
            {8'h00}, /* 0x4a62 */
            {8'h00}, /* 0x4a61 */
            {8'h00}, /* 0x4a60 */
            {8'h00}, /* 0x4a5f */
            {8'h00}, /* 0x4a5e */
            {8'h00}, /* 0x4a5d */
            {8'h00}, /* 0x4a5c */
            {8'h00}, /* 0x4a5b */
            {8'h00}, /* 0x4a5a */
            {8'h00}, /* 0x4a59 */
            {8'h00}, /* 0x4a58 */
            {8'h00}, /* 0x4a57 */
            {8'h00}, /* 0x4a56 */
            {8'h00}, /* 0x4a55 */
            {8'h00}, /* 0x4a54 */
            {8'h00}, /* 0x4a53 */
            {8'h00}, /* 0x4a52 */
            {8'h00}, /* 0x4a51 */
            {8'h00}, /* 0x4a50 */
            {8'h00}, /* 0x4a4f */
            {8'h00}, /* 0x4a4e */
            {8'h00}, /* 0x4a4d */
            {8'h00}, /* 0x4a4c */
            {8'h00}, /* 0x4a4b */
            {8'h00}, /* 0x4a4a */
            {8'h00}, /* 0x4a49 */
            {8'h00}, /* 0x4a48 */
            {8'h00}, /* 0x4a47 */
            {8'h00}, /* 0x4a46 */
            {8'h00}, /* 0x4a45 */
            {8'h00}, /* 0x4a44 */
            {8'h00}, /* 0x4a43 */
            {8'h00}, /* 0x4a42 */
            {8'h00}, /* 0x4a41 */
            {8'h00}, /* 0x4a40 */
            {8'h00}, /* 0x4a3f */
            {8'h00}, /* 0x4a3e */
            {8'h00}, /* 0x4a3d */
            {8'h00}, /* 0x4a3c */
            {8'h00}, /* 0x4a3b */
            {8'h00}, /* 0x4a3a */
            {8'h00}, /* 0x4a39 */
            {8'h00}, /* 0x4a38 */
            {8'h00}, /* 0x4a37 */
            {8'h00}, /* 0x4a36 */
            {8'h00}, /* 0x4a35 */
            {8'h00}, /* 0x4a34 */
            {8'h00}, /* 0x4a33 */
            {8'h00}, /* 0x4a32 */
            {8'h00}, /* 0x4a31 */
            {8'h00}, /* 0x4a30 */
            {8'h00}, /* 0x4a2f */
            {8'h00}, /* 0x4a2e */
            {8'h00}, /* 0x4a2d */
            {8'h00}, /* 0x4a2c */
            {8'h00}, /* 0x4a2b */
            {8'h00}, /* 0x4a2a */
            {8'h00}, /* 0x4a29 */
            {8'h00}, /* 0x4a28 */
            {8'h00}, /* 0x4a27 */
            {8'h00}, /* 0x4a26 */
            {8'h00}, /* 0x4a25 */
            {8'h00}, /* 0x4a24 */
            {8'h00}, /* 0x4a23 */
            {8'h00}, /* 0x4a22 */
            {8'h00}, /* 0x4a21 */
            {8'h00}, /* 0x4a20 */
            {8'h00}, /* 0x4a1f */
            {8'h00}, /* 0x4a1e */
            {8'h00}, /* 0x4a1d */
            {8'h00}, /* 0x4a1c */
            {8'h00}, /* 0x4a1b */
            {8'h00}, /* 0x4a1a */
            {8'h00}, /* 0x4a19 */
            {8'h00}, /* 0x4a18 */
            {8'h00}, /* 0x4a17 */
            {8'h00}, /* 0x4a16 */
            {8'h00}, /* 0x4a15 */
            {8'h00}, /* 0x4a14 */
            {8'h00}, /* 0x4a13 */
            {8'h00}, /* 0x4a12 */
            {8'h00}, /* 0x4a11 */
            {8'h00}, /* 0x4a10 */
            {8'h00}, /* 0x4a0f */
            {8'h00}, /* 0x4a0e */
            {8'h00}, /* 0x4a0d */
            {8'h00}, /* 0x4a0c */
            {8'h00}, /* 0x4a0b */
            {8'h00}, /* 0x4a0a */
            {8'h00}, /* 0x4a09 */
            {8'h00}, /* 0x4a08 */
            {8'h00}, /* 0x4a07 */
            {8'h00}, /* 0x4a06 */
            {8'h00}, /* 0x4a05 */
            {8'h00}, /* 0x4a04 */
            {8'h00}, /* 0x4a03 */
            {8'h00}, /* 0x4a02 */
            {8'h00}, /* 0x4a01 */
            {8'h00}, /* 0x4a00 */
            {8'h00}, /* 0x49ff */
            {8'h00}, /* 0x49fe */
            {8'h00}, /* 0x49fd */
            {8'h00}, /* 0x49fc */
            {8'h00}, /* 0x49fb */
            {8'h00}, /* 0x49fa */
            {8'h00}, /* 0x49f9 */
            {8'h00}, /* 0x49f8 */
            {8'h00}, /* 0x49f7 */
            {8'h00}, /* 0x49f6 */
            {8'h00}, /* 0x49f5 */
            {8'h00}, /* 0x49f4 */
            {8'h00}, /* 0x49f3 */
            {8'h00}, /* 0x49f2 */
            {8'h00}, /* 0x49f1 */
            {8'h00}, /* 0x49f0 */
            {8'h00}, /* 0x49ef */
            {8'h00}, /* 0x49ee */
            {8'h00}, /* 0x49ed */
            {8'h00}, /* 0x49ec */
            {8'h00}, /* 0x49eb */
            {8'h00}, /* 0x49ea */
            {8'h00}, /* 0x49e9 */
            {8'h00}, /* 0x49e8 */
            {8'h00}, /* 0x49e7 */
            {8'h00}, /* 0x49e6 */
            {8'h00}, /* 0x49e5 */
            {8'h00}, /* 0x49e4 */
            {8'h00}, /* 0x49e3 */
            {8'h00}, /* 0x49e2 */
            {8'h00}, /* 0x49e1 */
            {8'h00}, /* 0x49e0 */
            {8'h00}, /* 0x49df */
            {8'h00}, /* 0x49de */
            {8'h00}, /* 0x49dd */
            {8'h00}, /* 0x49dc */
            {8'h00}, /* 0x49db */
            {8'h00}, /* 0x49da */
            {8'h00}, /* 0x49d9 */
            {8'h00}, /* 0x49d8 */
            {8'h00}, /* 0x49d7 */
            {8'h00}, /* 0x49d6 */
            {8'h00}, /* 0x49d5 */
            {8'h00}, /* 0x49d4 */
            {8'h00}, /* 0x49d3 */
            {8'h00}, /* 0x49d2 */
            {8'h00}, /* 0x49d1 */
            {8'h00}, /* 0x49d0 */
            {8'h00}, /* 0x49cf */
            {8'h00}, /* 0x49ce */
            {8'h00}, /* 0x49cd */
            {8'h00}, /* 0x49cc */
            {8'h00}, /* 0x49cb */
            {8'h00}, /* 0x49ca */
            {8'h00}, /* 0x49c9 */
            {8'h00}, /* 0x49c8 */
            {8'h00}, /* 0x49c7 */
            {8'h00}, /* 0x49c6 */
            {8'h00}, /* 0x49c5 */
            {8'h00}, /* 0x49c4 */
            {8'h00}, /* 0x49c3 */
            {8'h00}, /* 0x49c2 */
            {8'h00}, /* 0x49c1 */
            {8'h00}, /* 0x49c0 */
            {8'h00}, /* 0x49bf */
            {8'h00}, /* 0x49be */
            {8'h00}, /* 0x49bd */
            {8'h00}, /* 0x49bc */
            {8'h00}, /* 0x49bb */
            {8'h00}, /* 0x49ba */
            {8'h00}, /* 0x49b9 */
            {8'h00}, /* 0x49b8 */
            {8'h00}, /* 0x49b7 */
            {8'h00}, /* 0x49b6 */
            {8'h00}, /* 0x49b5 */
            {8'h00}, /* 0x49b4 */
            {8'h00}, /* 0x49b3 */
            {8'h00}, /* 0x49b2 */
            {8'h00}, /* 0x49b1 */
            {8'h00}, /* 0x49b0 */
            {8'h00}, /* 0x49af */
            {8'h00}, /* 0x49ae */
            {8'h00}, /* 0x49ad */
            {8'h00}, /* 0x49ac */
            {8'h00}, /* 0x49ab */
            {8'h00}, /* 0x49aa */
            {8'h00}, /* 0x49a9 */
            {8'h00}, /* 0x49a8 */
            {8'h00}, /* 0x49a7 */
            {8'h00}, /* 0x49a6 */
            {8'h00}, /* 0x49a5 */
            {8'h00}, /* 0x49a4 */
            {8'h00}, /* 0x49a3 */
            {8'h00}, /* 0x49a2 */
            {8'h00}, /* 0x49a1 */
            {8'h00}, /* 0x49a0 */
            {8'h00}, /* 0x499f */
            {8'h00}, /* 0x499e */
            {8'h00}, /* 0x499d */
            {8'h00}, /* 0x499c */
            {8'h00}, /* 0x499b */
            {8'h00}, /* 0x499a */
            {8'h00}, /* 0x4999 */
            {8'h00}, /* 0x4998 */
            {8'h00}, /* 0x4997 */
            {8'h00}, /* 0x4996 */
            {8'h00}, /* 0x4995 */
            {8'h00}, /* 0x4994 */
            {8'h00}, /* 0x4993 */
            {8'h00}, /* 0x4992 */
            {8'h00}, /* 0x4991 */
            {8'h00}, /* 0x4990 */
            {8'h00}, /* 0x498f */
            {8'h00}, /* 0x498e */
            {8'h00}, /* 0x498d */
            {8'h00}, /* 0x498c */
            {8'h00}, /* 0x498b */
            {8'h00}, /* 0x498a */
            {8'h00}, /* 0x4989 */
            {8'h00}, /* 0x4988 */
            {8'h00}, /* 0x4987 */
            {8'h00}, /* 0x4986 */
            {8'h00}, /* 0x4985 */
            {8'h00}, /* 0x4984 */
            {8'h00}, /* 0x4983 */
            {8'h00}, /* 0x4982 */
            {8'h00}, /* 0x4981 */
            {8'h00}, /* 0x4980 */
            {8'h00}, /* 0x497f */
            {8'h00}, /* 0x497e */
            {8'h00}, /* 0x497d */
            {8'h00}, /* 0x497c */
            {8'h00}, /* 0x497b */
            {8'h00}, /* 0x497a */
            {8'h00}, /* 0x4979 */
            {8'h00}, /* 0x4978 */
            {8'h00}, /* 0x4977 */
            {8'h00}, /* 0x4976 */
            {8'h00}, /* 0x4975 */
            {8'h00}, /* 0x4974 */
            {8'h00}, /* 0x4973 */
            {8'h00}, /* 0x4972 */
            {8'h00}, /* 0x4971 */
            {8'h00}, /* 0x4970 */
            {8'h00}, /* 0x496f */
            {8'h00}, /* 0x496e */
            {8'h00}, /* 0x496d */
            {8'h00}, /* 0x496c */
            {8'h00}, /* 0x496b */
            {8'h00}, /* 0x496a */
            {8'h00}, /* 0x4969 */
            {8'h00}, /* 0x4968 */
            {8'h00}, /* 0x4967 */
            {8'h00}, /* 0x4966 */
            {8'h00}, /* 0x4965 */
            {8'h00}, /* 0x4964 */
            {8'h00}, /* 0x4963 */
            {8'h00}, /* 0x4962 */
            {8'h00}, /* 0x4961 */
            {8'h00}, /* 0x4960 */
            {8'h00}, /* 0x495f */
            {8'h00}, /* 0x495e */
            {8'h00}, /* 0x495d */
            {8'h00}, /* 0x495c */
            {8'h00}, /* 0x495b */
            {8'h00}, /* 0x495a */
            {8'h00}, /* 0x4959 */
            {8'h00}, /* 0x4958 */
            {8'h00}, /* 0x4957 */
            {8'h00}, /* 0x4956 */
            {8'h00}, /* 0x4955 */
            {8'h00}, /* 0x4954 */
            {8'h00}, /* 0x4953 */
            {8'h00}, /* 0x4952 */
            {8'h00}, /* 0x4951 */
            {8'h00}, /* 0x4950 */
            {8'h00}, /* 0x494f */
            {8'h00}, /* 0x494e */
            {8'h00}, /* 0x494d */
            {8'h00}, /* 0x494c */
            {8'h00}, /* 0x494b */
            {8'h00}, /* 0x494a */
            {8'h00}, /* 0x4949 */
            {8'h00}, /* 0x4948 */
            {8'h00}, /* 0x4947 */
            {8'h00}, /* 0x4946 */
            {8'h00}, /* 0x4945 */
            {8'h00}, /* 0x4944 */
            {8'h00}, /* 0x4943 */
            {8'h00}, /* 0x4942 */
            {8'h00}, /* 0x4941 */
            {8'h00}, /* 0x4940 */
            {8'h00}, /* 0x493f */
            {8'h00}, /* 0x493e */
            {8'h00}, /* 0x493d */
            {8'h00}, /* 0x493c */
            {8'h00}, /* 0x493b */
            {8'h00}, /* 0x493a */
            {8'h00}, /* 0x4939 */
            {8'h00}, /* 0x4938 */
            {8'h00}, /* 0x4937 */
            {8'h00}, /* 0x4936 */
            {8'h00}, /* 0x4935 */
            {8'h00}, /* 0x4934 */
            {8'h00}, /* 0x4933 */
            {8'h00}, /* 0x4932 */
            {8'h00}, /* 0x4931 */
            {8'h00}, /* 0x4930 */
            {8'h00}, /* 0x492f */
            {8'h00}, /* 0x492e */
            {8'h00}, /* 0x492d */
            {8'h00}, /* 0x492c */
            {8'h00}, /* 0x492b */
            {8'h00}, /* 0x492a */
            {8'h00}, /* 0x4929 */
            {8'h00}, /* 0x4928 */
            {8'h00}, /* 0x4927 */
            {8'h00}, /* 0x4926 */
            {8'h00}, /* 0x4925 */
            {8'h00}, /* 0x4924 */
            {8'h00}, /* 0x4923 */
            {8'h00}, /* 0x4922 */
            {8'h00}, /* 0x4921 */
            {8'h00}, /* 0x4920 */
            {8'h00}, /* 0x491f */
            {8'h00}, /* 0x491e */
            {8'h00}, /* 0x491d */
            {8'h00}, /* 0x491c */
            {8'h00}, /* 0x491b */
            {8'h00}, /* 0x491a */
            {8'h00}, /* 0x4919 */
            {8'h00}, /* 0x4918 */
            {8'h00}, /* 0x4917 */
            {8'h00}, /* 0x4916 */
            {8'h00}, /* 0x4915 */
            {8'h00}, /* 0x4914 */
            {8'h00}, /* 0x4913 */
            {8'h00}, /* 0x4912 */
            {8'h00}, /* 0x4911 */
            {8'h00}, /* 0x4910 */
            {8'h00}, /* 0x490f */
            {8'h00}, /* 0x490e */
            {8'h00}, /* 0x490d */
            {8'h00}, /* 0x490c */
            {8'h00}, /* 0x490b */
            {8'h00}, /* 0x490a */
            {8'h00}, /* 0x4909 */
            {8'h00}, /* 0x4908 */
            {8'h00}, /* 0x4907 */
            {8'h00}, /* 0x4906 */
            {8'h00}, /* 0x4905 */
            {8'h00}, /* 0x4904 */
            {8'h00}, /* 0x4903 */
            {8'h00}, /* 0x4902 */
            {8'h00}, /* 0x4901 */
            {8'h00}, /* 0x4900 */
            {8'h00}, /* 0x48ff */
            {8'h00}, /* 0x48fe */
            {8'h00}, /* 0x48fd */
            {8'h00}, /* 0x48fc */
            {8'h00}, /* 0x48fb */
            {8'h00}, /* 0x48fa */
            {8'h00}, /* 0x48f9 */
            {8'h00}, /* 0x48f8 */
            {8'h00}, /* 0x48f7 */
            {8'h00}, /* 0x48f6 */
            {8'h00}, /* 0x48f5 */
            {8'h00}, /* 0x48f4 */
            {8'h00}, /* 0x48f3 */
            {8'h00}, /* 0x48f2 */
            {8'h00}, /* 0x48f1 */
            {8'h00}, /* 0x48f0 */
            {8'h00}, /* 0x48ef */
            {8'h00}, /* 0x48ee */
            {8'h00}, /* 0x48ed */
            {8'h00}, /* 0x48ec */
            {8'h00}, /* 0x48eb */
            {8'h00}, /* 0x48ea */
            {8'h00}, /* 0x48e9 */
            {8'h00}, /* 0x48e8 */
            {8'h00}, /* 0x48e7 */
            {8'h00}, /* 0x48e6 */
            {8'h00}, /* 0x48e5 */
            {8'h00}, /* 0x48e4 */
            {8'h00}, /* 0x48e3 */
            {8'h00}, /* 0x48e2 */
            {8'h00}, /* 0x48e1 */
            {8'h00}, /* 0x48e0 */
            {8'h00}, /* 0x48df */
            {8'h00}, /* 0x48de */
            {8'h00}, /* 0x48dd */
            {8'h00}, /* 0x48dc */
            {8'h00}, /* 0x48db */
            {8'h00}, /* 0x48da */
            {8'h00}, /* 0x48d9 */
            {8'h00}, /* 0x48d8 */
            {8'h00}, /* 0x48d7 */
            {8'h00}, /* 0x48d6 */
            {8'h00}, /* 0x48d5 */
            {8'h00}, /* 0x48d4 */
            {8'h00}, /* 0x48d3 */
            {8'h00}, /* 0x48d2 */
            {8'h00}, /* 0x48d1 */
            {8'h00}, /* 0x48d0 */
            {8'h00}, /* 0x48cf */
            {8'h00}, /* 0x48ce */
            {8'h00}, /* 0x48cd */
            {8'h00}, /* 0x48cc */
            {8'h00}, /* 0x48cb */
            {8'h00}, /* 0x48ca */
            {8'h00}, /* 0x48c9 */
            {8'h00}, /* 0x48c8 */
            {8'h00}, /* 0x48c7 */
            {8'h00}, /* 0x48c6 */
            {8'h00}, /* 0x48c5 */
            {8'h00}, /* 0x48c4 */
            {8'h00}, /* 0x48c3 */
            {8'h00}, /* 0x48c2 */
            {8'h00}, /* 0x48c1 */
            {8'h00}, /* 0x48c0 */
            {8'h00}, /* 0x48bf */
            {8'h00}, /* 0x48be */
            {8'h00}, /* 0x48bd */
            {8'h00}, /* 0x48bc */
            {8'h00}, /* 0x48bb */
            {8'h00}, /* 0x48ba */
            {8'h00}, /* 0x48b9 */
            {8'h00}, /* 0x48b8 */
            {8'h00}, /* 0x48b7 */
            {8'h00}, /* 0x48b6 */
            {8'h00}, /* 0x48b5 */
            {8'h00}, /* 0x48b4 */
            {8'h00}, /* 0x48b3 */
            {8'h00}, /* 0x48b2 */
            {8'h00}, /* 0x48b1 */
            {8'h00}, /* 0x48b0 */
            {8'h00}, /* 0x48af */
            {8'h00}, /* 0x48ae */
            {8'h00}, /* 0x48ad */
            {8'h00}, /* 0x48ac */
            {8'h00}, /* 0x48ab */
            {8'h00}, /* 0x48aa */
            {8'h00}, /* 0x48a9 */
            {8'h00}, /* 0x48a8 */
            {8'h00}, /* 0x48a7 */
            {8'h00}, /* 0x48a6 */
            {8'h00}, /* 0x48a5 */
            {8'h00}, /* 0x48a4 */
            {8'h00}, /* 0x48a3 */
            {8'h00}, /* 0x48a2 */
            {8'h00}, /* 0x48a1 */
            {8'h00}, /* 0x48a0 */
            {8'h00}, /* 0x489f */
            {8'h00}, /* 0x489e */
            {8'h00}, /* 0x489d */
            {8'h00}, /* 0x489c */
            {8'h00}, /* 0x489b */
            {8'h00}, /* 0x489a */
            {8'h00}, /* 0x4899 */
            {8'h00}, /* 0x4898 */
            {8'h00}, /* 0x4897 */
            {8'h00}, /* 0x4896 */
            {8'h00}, /* 0x4895 */
            {8'h00}, /* 0x4894 */
            {8'h00}, /* 0x4893 */
            {8'h00}, /* 0x4892 */
            {8'h00}, /* 0x4891 */
            {8'h00}, /* 0x4890 */
            {8'h00}, /* 0x488f */
            {8'h00}, /* 0x488e */
            {8'h00}, /* 0x488d */
            {8'h00}, /* 0x488c */
            {8'h00}, /* 0x488b */
            {8'h00}, /* 0x488a */
            {8'h00}, /* 0x4889 */
            {8'h00}, /* 0x4888 */
            {8'h00}, /* 0x4887 */
            {8'h00}, /* 0x4886 */
            {8'h00}, /* 0x4885 */
            {8'h00}, /* 0x4884 */
            {8'h00}, /* 0x4883 */
            {8'h00}, /* 0x4882 */
            {8'h00}, /* 0x4881 */
            {8'h00}, /* 0x4880 */
            {8'h00}, /* 0x487f */
            {8'h00}, /* 0x487e */
            {8'h00}, /* 0x487d */
            {8'h00}, /* 0x487c */
            {8'h00}, /* 0x487b */
            {8'h00}, /* 0x487a */
            {8'h00}, /* 0x4879 */
            {8'h00}, /* 0x4878 */
            {8'h00}, /* 0x4877 */
            {8'h00}, /* 0x4876 */
            {8'h00}, /* 0x4875 */
            {8'h00}, /* 0x4874 */
            {8'h00}, /* 0x4873 */
            {8'h00}, /* 0x4872 */
            {8'h00}, /* 0x4871 */
            {8'h00}, /* 0x4870 */
            {8'h00}, /* 0x486f */
            {8'h00}, /* 0x486e */
            {8'h00}, /* 0x486d */
            {8'h00}, /* 0x486c */
            {8'h00}, /* 0x486b */
            {8'h00}, /* 0x486a */
            {8'h00}, /* 0x4869 */
            {8'h00}, /* 0x4868 */
            {8'h00}, /* 0x4867 */
            {8'h00}, /* 0x4866 */
            {8'h00}, /* 0x4865 */
            {8'h00}, /* 0x4864 */
            {8'h00}, /* 0x4863 */
            {8'h00}, /* 0x4862 */
            {8'h00}, /* 0x4861 */
            {8'h00}, /* 0x4860 */
            {8'h00}, /* 0x485f */
            {8'h00}, /* 0x485e */
            {8'h00}, /* 0x485d */
            {8'h00}, /* 0x485c */
            {8'h00}, /* 0x485b */
            {8'h00}, /* 0x485a */
            {8'h00}, /* 0x4859 */
            {8'h00}, /* 0x4858 */
            {8'h00}, /* 0x4857 */
            {8'h00}, /* 0x4856 */
            {8'h00}, /* 0x4855 */
            {8'h00}, /* 0x4854 */
            {8'h00}, /* 0x4853 */
            {8'h00}, /* 0x4852 */
            {8'h00}, /* 0x4851 */
            {8'h00}, /* 0x4850 */
            {8'h00}, /* 0x484f */
            {8'h00}, /* 0x484e */
            {8'h00}, /* 0x484d */
            {8'h00}, /* 0x484c */
            {8'h00}, /* 0x484b */
            {8'h00}, /* 0x484a */
            {8'h00}, /* 0x4849 */
            {8'h00}, /* 0x4848 */
            {8'h00}, /* 0x4847 */
            {8'h00}, /* 0x4846 */
            {8'h00}, /* 0x4845 */
            {8'h00}, /* 0x4844 */
            {8'h00}, /* 0x4843 */
            {8'h00}, /* 0x4842 */
            {8'h00}, /* 0x4841 */
            {8'h00}, /* 0x4840 */
            {8'h00}, /* 0x483f */
            {8'h00}, /* 0x483e */
            {8'h00}, /* 0x483d */
            {8'h00}, /* 0x483c */
            {8'h00}, /* 0x483b */
            {8'h00}, /* 0x483a */
            {8'h00}, /* 0x4839 */
            {8'h00}, /* 0x4838 */
            {8'h00}, /* 0x4837 */
            {8'h00}, /* 0x4836 */
            {8'h00}, /* 0x4835 */
            {8'h00}, /* 0x4834 */
            {8'h00}, /* 0x4833 */
            {8'h00}, /* 0x4832 */
            {8'h00}, /* 0x4831 */
            {8'h00}, /* 0x4830 */
            {8'h00}, /* 0x482f */
            {8'h00}, /* 0x482e */
            {8'h00}, /* 0x482d */
            {8'h00}, /* 0x482c */
            {8'h00}, /* 0x482b */
            {8'h00}, /* 0x482a */
            {8'h00}, /* 0x4829 */
            {8'h00}, /* 0x4828 */
            {8'h00}, /* 0x4827 */
            {8'h00}, /* 0x4826 */
            {8'h00}, /* 0x4825 */
            {8'h00}, /* 0x4824 */
            {8'h00}, /* 0x4823 */
            {8'h00}, /* 0x4822 */
            {8'h00}, /* 0x4821 */
            {8'h00}, /* 0x4820 */
            {8'h00}, /* 0x481f */
            {8'h00}, /* 0x481e */
            {8'h00}, /* 0x481d */
            {8'h00}, /* 0x481c */
            {8'h00}, /* 0x481b */
            {8'h00}, /* 0x481a */
            {8'h00}, /* 0x4819 */
            {8'h00}, /* 0x4818 */
            {8'h00}, /* 0x4817 */
            {8'h00}, /* 0x4816 */
            {8'h00}, /* 0x4815 */
            {8'h00}, /* 0x4814 */
            {8'h00}, /* 0x4813 */
            {8'h00}, /* 0x4812 */
            {8'h00}, /* 0x4811 */
            {8'h00}, /* 0x4810 */
            {8'h00}, /* 0x480f */
            {8'h00}, /* 0x480e */
            {8'h00}, /* 0x480d */
            {8'h00}, /* 0x480c */
            {8'h00}, /* 0x480b */
            {8'h00}, /* 0x480a */
            {8'h00}, /* 0x4809 */
            {8'h00}, /* 0x4808 */
            {8'h00}, /* 0x4807 */
            {8'h00}, /* 0x4806 */
            {8'h00}, /* 0x4805 */
            {8'h00}, /* 0x4804 */
            {8'h00}, /* 0x4803 */
            {8'h00}, /* 0x4802 */
            {8'h00}, /* 0x4801 */
            {8'h00}, /* 0x4800 */
            {8'h00}, /* 0x47ff */
            {8'h00}, /* 0x47fe */
            {8'h00}, /* 0x47fd */
            {8'h00}, /* 0x47fc */
            {8'h00}, /* 0x47fb */
            {8'h00}, /* 0x47fa */
            {8'h00}, /* 0x47f9 */
            {8'h00}, /* 0x47f8 */
            {8'h00}, /* 0x47f7 */
            {8'h00}, /* 0x47f6 */
            {8'h00}, /* 0x47f5 */
            {8'h00}, /* 0x47f4 */
            {8'h00}, /* 0x47f3 */
            {8'h00}, /* 0x47f2 */
            {8'h00}, /* 0x47f1 */
            {8'h00}, /* 0x47f0 */
            {8'h00}, /* 0x47ef */
            {8'h00}, /* 0x47ee */
            {8'h00}, /* 0x47ed */
            {8'h00}, /* 0x47ec */
            {8'h00}, /* 0x47eb */
            {8'h00}, /* 0x47ea */
            {8'h00}, /* 0x47e9 */
            {8'h00}, /* 0x47e8 */
            {8'h00}, /* 0x47e7 */
            {8'h00}, /* 0x47e6 */
            {8'h00}, /* 0x47e5 */
            {8'h00}, /* 0x47e4 */
            {8'h00}, /* 0x47e3 */
            {8'h00}, /* 0x47e2 */
            {8'h00}, /* 0x47e1 */
            {8'h00}, /* 0x47e0 */
            {8'h00}, /* 0x47df */
            {8'h00}, /* 0x47de */
            {8'h00}, /* 0x47dd */
            {8'h00}, /* 0x47dc */
            {8'h00}, /* 0x47db */
            {8'h00}, /* 0x47da */
            {8'h00}, /* 0x47d9 */
            {8'h00}, /* 0x47d8 */
            {8'h00}, /* 0x47d7 */
            {8'h00}, /* 0x47d6 */
            {8'h00}, /* 0x47d5 */
            {8'h00}, /* 0x47d4 */
            {8'h00}, /* 0x47d3 */
            {8'h00}, /* 0x47d2 */
            {8'h00}, /* 0x47d1 */
            {8'h00}, /* 0x47d0 */
            {8'h00}, /* 0x47cf */
            {8'h00}, /* 0x47ce */
            {8'h00}, /* 0x47cd */
            {8'h00}, /* 0x47cc */
            {8'h00}, /* 0x47cb */
            {8'h00}, /* 0x47ca */
            {8'h00}, /* 0x47c9 */
            {8'h00}, /* 0x47c8 */
            {8'h00}, /* 0x47c7 */
            {8'h00}, /* 0x47c6 */
            {8'h00}, /* 0x47c5 */
            {8'h00}, /* 0x47c4 */
            {8'h00}, /* 0x47c3 */
            {8'h00}, /* 0x47c2 */
            {8'h00}, /* 0x47c1 */
            {8'h00}, /* 0x47c0 */
            {8'h00}, /* 0x47bf */
            {8'h00}, /* 0x47be */
            {8'h00}, /* 0x47bd */
            {8'h00}, /* 0x47bc */
            {8'h00}, /* 0x47bb */
            {8'h00}, /* 0x47ba */
            {8'h00}, /* 0x47b9 */
            {8'h00}, /* 0x47b8 */
            {8'h00}, /* 0x47b7 */
            {8'h00}, /* 0x47b6 */
            {8'h00}, /* 0x47b5 */
            {8'h00}, /* 0x47b4 */
            {8'h00}, /* 0x47b3 */
            {8'h00}, /* 0x47b2 */
            {8'h00}, /* 0x47b1 */
            {8'h00}, /* 0x47b0 */
            {8'h00}, /* 0x47af */
            {8'h00}, /* 0x47ae */
            {8'h00}, /* 0x47ad */
            {8'h00}, /* 0x47ac */
            {8'h00}, /* 0x47ab */
            {8'h00}, /* 0x47aa */
            {8'h00}, /* 0x47a9 */
            {8'h00}, /* 0x47a8 */
            {8'h00}, /* 0x47a7 */
            {8'h00}, /* 0x47a6 */
            {8'h00}, /* 0x47a5 */
            {8'h00}, /* 0x47a4 */
            {8'h00}, /* 0x47a3 */
            {8'h00}, /* 0x47a2 */
            {8'h00}, /* 0x47a1 */
            {8'h00}, /* 0x47a0 */
            {8'h00}, /* 0x479f */
            {8'h00}, /* 0x479e */
            {8'h00}, /* 0x479d */
            {8'h00}, /* 0x479c */
            {8'h00}, /* 0x479b */
            {8'h00}, /* 0x479a */
            {8'h00}, /* 0x4799 */
            {8'h00}, /* 0x4798 */
            {8'h00}, /* 0x4797 */
            {8'h00}, /* 0x4796 */
            {8'h00}, /* 0x4795 */
            {8'h00}, /* 0x4794 */
            {8'h00}, /* 0x4793 */
            {8'h00}, /* 0x4792 */
            {8'h00}, /* 0x4791 */
            {8'h00}, /* 0x4790 */
            {8'h00}, /* 0x478f */
            {8'h00}, /* 0x478e */
            {8'h00}, /* 0x478d */
            {8'h00}, /* 0x478c */
            {8'h00}, /* 0x478b */
            {8'h00}, /* 0x478a */
            {8'h00}, /* 0x4789 */
            {8'h00}, /* 0x4788 */
            {8'h00}, /* 0x4787 */
            {8'h00}, /* 0x4786 */
            {8'h00}, /* 0x4785 */
            {8'h00}, /* 0x4784 */
            {8'h00}, /* 0x4783 */
            {8'h00}, /* 0x4782 */
            {8'h00}, /* 0x4781 */
            {8'h00}, /* 0x4780 */
            {8'h00}, /* 0x477f */
            {8'h00}, /* 0x477e */
            {8'h00}, /* 0x477d */
            {8'h00}, /* 0x477c */
            {8'h00}, /* 0x477b */
            {8'h00}, /* 0x477a */
            {8'h00}, /* 0x4779 */
            {8'h00}, /* 0x4778 */
            {8'h00}, /* 0x4777 */
            {8'h00}, /* 0x4776 */
            {8'h00}, /* 0x4775 */
            {8'h00}, /* 0x4774 */
            {8'h00}, /* 0x4773 */
            {8'h00}, /* 0x4772 */
            {8'h00}, /* 0x4771 */
            {8'h00}, /* 0x4770 */
            {8'h00}, /* 0x476f */
            {8'h00}, /* 0x476e */
            {8'h00}, /* 0x476d */
            {8'h00}, /* 0x476c */
            {8'h00}, /* 0x476b */
            {8'h00}, /* 0x476a */
            {8'h00}, /* 0x4769 */
            {8'h00}, /* 0x4768 */
            {8'h00}, /* 0x4767 */
            {8'h00}, /* 0x4766 */
            {8'h00}, /* 0x4765 */
            {8'h00}, /* 0x4764 */
            {8'h00}, /* 0x4763 */
            {8'h00}, /* 0x4762 */
            {8'h00}, /* 0x4761 */
            {8'h00}, /* 0x4760 */
            {8'h00}, /* 0x475f */
            {8'h00}, /* 0x475e */
            {8'h00}, /* 0x475d */
            {8'h00}, /* 0x475c */
            {8'h00}, /* 0x475b */
            {8'h00}, /* 0x475a */
            {8'h00}, /* 0x4759 */
            {8'h00}, /* 0x4758 */
            {8'h00}, /* 0x4757 */
            {8'h00}, /* 0x4756 */
            {8'h00}, /* 0x4755 */
            {8'h00}, /* 0x4754 */
            {8'h00}, /* 0x4753 */
            {8'h00}, /* 0x4752 */
            {8'h00}, /* 0x4751 */
            {8'h00}, /* 0x4750 */
            {8'h00}, /* 0x474f */
            {8'h00}, /* 0x474e */
            {8'h00}, /* 0x474d */
            {8'h00}, /* 0x474c */
            {8'h00}, /* 0x474b */
            {8'h00}, /* 0x474a */
            {8'h00}, /* 0x4749 */
            {8'h00}, /* 0x4748 */
            {8'h00}, /* 0x4747 */
            {8'h00}, /* 0x4746 */
            {8'h00}, /* 0x4745 */
            {8'h00}, /* 0x4744 */
            {8'h00}, /* 0x4743 */
            {8'h00}, /* 0x4742 */
            {8'h00}, /* 0x4741 */
            {8'h00}, /* 0x4740 */
            {8'h00}, /* 0x473f */
            {8'h00}, /* 0x473e */
            {8'h00}, /* 0x473d */
            {8'h00}, /* 0x473c */
            {8'h00}, /* 0x473b */
            {8'h00}, /* 0x473a */
            {8'h00}, /* 0x4739 */
            {8'h00}, /* 0x4738 */
            {8'h00}, /* 0x4737 */
            {8'h00}, /* 0x4736 */
            {8'h00}, /* 0x4735 */
            {8'h00}, /* 0x4734 */
            {8'h00}, /* 0x4733 */
            {8'h00}, /* 0x4732 */
            {8'h00}, /* 0x4731 */
            {8'h00}, /* 0x4730 */
            {8'h00}, /* 0x472f */
            {8'h00}, /* 0x472e */
            {8'h00}, /* 0x472d */
            {8'h00}, /* 0x472c */
            {8'h00}, /* 0x472b */
            {8'h00}, /* 0x472a */
            {8'h00}, /* 0x4729 */
            {8'h00}, /* 0x4728 */
            {8'h00}, /* 0x4727 */
            {8'h00}, /* 0x4726 */
            {8'h00}, /* 0x4725 */
            {8'h00}, /* 0x4724 */
            {8'h00}, /* 0x4723 */
            {8'h00}, /* 0x4722 */
            {8'h00}, /* 0x4721 */
            {8'h00}, /* 0x4720 */
            {8'h00}, /* 0x471f */
            {8'h00}, /* 0x471e */
            {8'h00}, /* 0x471d */
            {8'h00}, /* 0x471c */
            {8'h00}, /* 0x471b */
            {8'h00}, /* 0x471a */
            {8'h00}, /* 0x4719 */
            {8'h00}, /* 0x4718 */
            {8'h00}, /* 0x4717 */
            {8'h00}, /* 0x4716 */
            {8'h00}, /* 0x4715 */
            {8'h00}, /* 0x4714 */
            {8'h00}, /* 0x4713 */
            {8'h00}, /* 0x4712 */
            {8'h00}, /* 0x4711 */
            {8'h00}, /* 0x4710 */
            {8'h00}, /* 0x470f */
            {8'h00}, /* 0x470e */
            {8'h00}, /* 0x470d */
            {8'h00}, /* 0x470c */
            {8'h00}, /* 0x470b */
            {8'h00}, /* 0x470a */
            {8'h00}, /* 0x4709 */
            {8'h00}, /* 0x4708 */
            {8'h00}, /* 0x4707 */
            {8'h00}, /* 0x4706 */
            {8'h00}, /* 0x4705 */
            {8'h00}, /* 0x4704 */
            {8'h00}, /* 0x4703 */
            {8'h00}, /* 0x4702 */
            {8'h00}, /* 0x4701 */
            {8'h00}, /* 0x4700 */
            {8'h00}, /* 0x46ff */
            {8'h00}, /* 0x46fe */
            {8'h00}, /* 0x46fd */
            {8'h00}, /* 0x46fc */
            {8'h00}, /* 0x46fb */
            {8'h00}, /* 0x46fa */
            {8'h00}, /* 0x46f9 */
            {8'h00}, /* 0x46f8 */
            {8'h00}, /* 0x46f7 */
            {8'h00}, /* 0x46f6 */
            {8'h00}, /* 0x46f5 */
            {8'h00}, /* 0x46f4 */
            {8'h00}, /* 0x46f3 */
            {8'h00}, /* 0x46f2 */
            {8'h00}, /* 0x46f1 */
            {8'h00}, /* 0x46f0 */
            {8'h00}, /* 0x46ef */
            {8'h00}, /* 0x46ee */
            {8'h00}, /* 0x46ed */
            {8'h00}, /* 0x46ec */
            {8'h00}, /* 0x46eb */
            {8'h00}, /* 0x46ea */
            {8'h00}, /* 0x46e9 */
            {8'h00}, /* 0x46e8 */
            {8'h00}, /* 0x46e7 */
            {8'h00}, /* 0x46e6 */
            {8'h00}, /* 0x46e5 */
            {8'h00}, /* 0x46e4 */
            {8'h00}, /* 0x46e3 */
            {8'h00}, /* 0x46e2 */
            {8'h00}, /* 0x46e1 */
            {8'h00}, /* 0x46e0 */
            {8'h00}, /* 0x46df */
            {8'h00}, /* 0x46de */
            {8'h00}, /* 0x46dd */
            {8'h00}, /* 0x46dc */
            {8'h00}, /* 0x46db */
            {8'h00}, /* 0x46da */
            {8'h00}, /* 0x46d9 */
            {8'h00}, /* 0x46d8 */
            {8'h00}, /* 0x46d7 */
            {8'h00}, /* 0x46d6 */
            {8'h00}, /* 0x46d5 */
            {8'h00}, /* 0x46d4 */
            {8'h00}, /* 0x46d3 */
            {8'h00}, /* 0x46d2 */
            {8'h00}, /* 0x46d1 */
            {8'h00}, /* 0x46d0 */
            {8'h00}, /* 0x46cf */
            {8'h00}, /* 0x46ce */
            {8'h00}, /* 0x46cd */
            {8'h00}, /* 0x46cc */
            {8'h00}, /* 0x46cb */
            {8'h00}, /* 0x46ca */
            {8'h00}, /* 0x46c9 */
            {8'h00}, /* 0x46c8 */
            {8'h00}, /* 0x46c7 */
            {8'h00}, /* 0x46c6 */
            {8'h00}, /* 0x46c5 */
            {8'h00}, /* 0x46c4 */
            {8'h00}, /* 0x46c3 */
            {8'h00}, /* 0x46c2 */
            {8'h00}, /* 0x46c1 */
            {8'h00}, /* 0x46c0 */
            {8'h00}, /* 0x46bf */
            {8'h00}, /* 0x46be */
            {8'h00}, /* 0x46bd */
            {8'h00}, /* 0x46bc */
            {8'h00}, /* 0x46bb */
            {8'h00}, /* 0x46ba */
            {8'h00}, /* 0x46b9 */
            {8'h00}, /* 0x46b8 */
            {8'h00}, /* 0x46b7 */
            {8'h00}, /* 0x46b6 */
            {8'h00}, /* 0x46b5 */
            {8'h00}, /* 0x46b4 */
            {8'h00}, /* 0x46b3 */
            {8'h00}, /* 0x46b2 */
            {8'h00}, /* 0x46b1 */
            {8'h00}, /* 0x46b0 */
            {8'h00}, /* 0x46af */
            {8'h00}, /* 0x46ae */
            {8'h00}, /* 0x46ad */
            {8'h00}, /* 0x46ac */
            {8'h00}, /* 0x46ab */
            {8'h00}, /* 0x46aa */
            {8'h00}, /* 0x46a9 */
            {8'h00}, /* 0x46a8 */
            {8'h00}, /* 0x46a7 */
            {8'h00}, /* 0x46a6 */
            {8'h00}, /* 0x46a5 */
            {8'h00}, /* 0x46a4 */
            {8'h00}, /* 0x46a3 */
            {8'h00}, /* 0x46a2 */
            {8'h00}, /* 0x46a1 */
            {8'h00}, /* 0x46a0 */
            {8'h00}, /* 0x469f */
            {8'h00}, /* 0x469e */
            {8'h00}, /* 0x469d */
            {8'h00}, /* 0x469c */
            {8'h00}, /* 0x469b */
            {8'h00}, /* 0x469a */
            {8'h00}, /* 0x4699 */
            {8'h00}, /* 0x4698 */
            {8'h00}, /* 0x4697 */
            {8'h00}, /* 0x4696 */
            {8'h00}, /* 0x4695 */
            {8'h00}, /* 0x4694 */
            {8'h00}, /* 0x4693 */
            {8'h00}, /* 0x4692 */
            {8'h00}, /* 0x4691 */
            {8'h00}, /* 0x4690 */
            {8'h00}, /* 0x468f */
            {8'h00}, /* 0x468e */
            {8'h00}, /* 0x468d */
            {8'h00}, /* 0x468c */
            {8'h00}, /* 0x468b */
            {8'h00}, /* 0x468a */
            {8'h00}, /* 0x4689 */
            {8'h00}, /* 0x4688 */
            {8'h00}, /* 0x4687 */
            {8'h00}, /* 0x4686 */
            {8'h00}, /* 0x4685 */
            {8'h00}, /* 0x4684 */
            {8'h00}, /* 0x4683 */
            {8'h00}, /* 0x4682 */
            {8'h00}, /* 0x4681 */
            {8'h00}, /* 0x4680 */
            {8'h00}, /* 0x467f */
            {8'h00}, /* 0x467e */
            {8'h00}, /* 0x467d */
            {8'h00}, /* 0x467c */
            {8'h00}, /* 0x467b */
            {8'h00}, /* 0x467a */
            {8'h00}, /* 0x4679 */
            {8'h00}, /* 0x4678 */
            {8'h00}, /* 0x4677 */
            {8'h00}, /* 0x4676 */
            {8'h00}, /* 0x4675 */
            {8'h00}, /* 0x4674 */
            {8'h00}, /* 0x4673 */
            {8'h00}, /* 0x4672 */
            {8'h00}, /* 0x4671 */
            {8'h00}, /* 0x4670 */
            {8'h00}, /* 0x466f */
            {8'h00}, /* 0x466e */
            {8'h00}, /* 0x466d */
            {8'h00}, /* 0x466c */
            {8'h00}, /* 0x466b */
            {8'h00}, /* 0x466a */
            {8'h00}, /* 0x4669 */
            {8'h00}, /* 0x4668 */
            {8'h00}, /* 0x4667 */
            {8'h00}, /* 0x4666 */
            {8'h00}, /* 0x4665 */
            {8'h00}, /* 0x4664 */
            {8'h00}, /* 0x4663 */
            {8'h00}, /* 0x4662 */
            {8'h00}, /* 0x4661 */
            {8'h00}, /* 0x4660 */
            {8'h00}, /* 0x465f */
            {8'h00}, /* 0x465e */
            {8'h00}, /* 0x465d */
            {8'h00}, /* 0x465c */
            {8'h00}, /* 0x465b */
            {8'h00}, /* 0x465a */
            {8'h00}, /* 0x4659 */
            {8'h00}, /* 0x4658 */
            {8'h00}, /* 0x4657 */
            {8'h00}, /* 0x4656 */
            {8'h00}, /* 0x4655 */
            {8'h00}, /* 0x4654 */
            {8'h00}, /* 0x4653 */
            {8'h00}, /* 0x4652 */
            {8'h00}, /* 0x4651 */
            {8'h00}, /* 0x4650 */
            {8'h00}, /* 0x464f */
            {8'h00}, /* 0x464e */
            {8'h00}, /* 0x464d */
            {8'h00}, /* 0x464c */
            {8'h00}, /* 0x464b */
            {8'h00}, /* 0x464a */
            {8'h00}, /* 0x4649 */
            {8'h00}, /* 0x4648 */
            {8'h00}, /* 0x4647 */
            {8'h00}, /* 0x4646 */
            {8'h00}, /* 0x4645 */
            {8'h00}, /* 0x4644 */
            {8'h00}, /* 0x4643 */
            {8'h00}, /* 0x4642 */
            {8'h00}, /* 0x4641 */
            {8'h00}, /* 0x4640 */
            {8'h00}, /* 0x463f */
            {8'h00}, /* 0x463e */
            {8'h00}, /* 0x463d */
            {8'h00}, /* 0x463c */
            {8'h00}, /* 0x463b */
            {8'h00}, /* 0x463a */
            {8'h00}, /* 0x4639 */
            {8'h00}, /* 0x4638 */
            {8'h00}, /* 0x4637 */
            {8'h00}, /* 0x4636 */
            {8'h00}, /* 0x4635 */
            {8'h00}, /* 0x4634 */
            {8'h00}, /* 0x4633 */
            {8'h00}, /* 0x4632 */
            {8'h00}, /* 0x4631 */
            {8'h00}, /* 0x4630 */
            {8'h00}, /* 0x462f */
            {8'h00}, /* 0x462e */
            {8'h00}, /* 0x462d */
            {8'h00}, /* 0x462c */
            {8'h00}, /* 0x462b */
            {8'h00}, /* 0x462a */
            {8'h00}, /* 0x4629 */
            {8'h00}, /* 0x4628 */
            {8'h00}, /* 0x4627 */
            {8'h00}, /* 0x4626 */
            {8'h00}, /* 0x4625 */
            {8'h00}, /* 0x4624 */
            {8'h00}, /* 0x4623 */
            {8'h00}, /* 0x4622 */
            {8'h00}, /* 0x4621 */
            {8'h00}, /* 0x4620 */
            {8'h00}, /* 0x461f */
            {8'h00}, /* 0x461e */
            {8'h00}, /* 0x461d */
            {8'h00}, /* 0x461c */
            {8'h00}, /* 0x461b */
            {8'h00}, /* 0x461a */
            {8'h00}, /* 0x4619 */
            {8'h00}, /* 0x4618 */
            {8'h00}, /* 0x4617 */
            {8'h00}, /* 0x4616 */
            {8'h00}, /* 0x4615 */
            {8'h00}, /* 0x4614 */
            {8'h00}, /* 0x4613 */
            {8'h00}, /* 0x4612 */
            {8'h00}, /* 0x4611 */
            {8'h00}, /* 0x4610 */
            {8'h00}, /* 0x460f */
            {8'h00}, /* 0x460e */
            {8'h00}, /* 0x460d */
            {8'h00}, /* 0x460c */
            {8'h00}, /* 0x460b */
            {8'h00}, /* 0x460a */
            {8'h00}, /* 0x4609 */
            {8'h00}, /* 0x4608 */
            {8'h00}, /* 0x4607 */
            {8'h00}, /* 0x4606 */
            {8'h00}, /* 0x4605 */
            {8'h00}, /* 0x4604 */
            {8'h00}, /* 0x4603 */
            {8'h00}, /* 0x4602 */
            {8'h00}, /* 0x4601 */
            {8'h00}, /* 0x4600 */
            {8'h00}, /* 0x45ff */
            {8'h00}, /* 0x45fe */
            {8'h00}, /* 0x45fd */
            {8'h00}, /* 0x45fc */
            {8'h00}, /* 0x45fb */
            {8'h00}, /* 0x45fa */
            {8'h00}, /* 0x45f9 */
            {8'h00}, /* 0x45f8 */
            {8'h00}, /* 0x45f7 */
            {8'h00}, /* 0x45f6 */
            {8'h00}, /* 0x45f5 */
            {8'h00}, /* 0x45f4 */
            {8'h00}, /* 0x45f3 */
            {8'h00}, /* 0x45f2 */
            {8'h00}, /* 0x45f1 */
            {8'h00}, /* 0x45f0 */
            {8'h00}, /* 0x45ef */
            {8'h00}, /* 0x45ee */
            {8'h00}, /* 0x45ed */
            {8'h00}, /* 0x45ec */
            {8'h00}, /* 0x45eb */
            {8'h00}, /* 0x45ea */
            {8'h00}, /* 0x45e9 */
            {8'h00}, /* 0x45e8 */
            {8'h00}, /* 0x45e7 */
            {8'h00}, /* 0x45e6 */
            {8'h00}, /* 0x45e5 */
            {8'h00}, /* 0x45e4 */
            {8'h00}, /* 0x45e3 */
            {8'h00}, /* 0x45e2 */
            {8'h00}, /* 0x45e1 */
            {8'h00}, /* 0x45e0 */
            {8'h00}, /* 0x45df */
            {8'h00}, /* 0x45de */
            {8'h00}, /* 0x45dd */
            {8'h00}, /* 0x45dc */
            {8'h00}, /* 0x45db */
            {8'h00}, /* 0x45da */
            {8'h00}, /* 0x45d9 */
            {8'h00}, /* 0x45d8 */
            {8'h00}, /* 0x45d7 */
            {8'h00}, /* 0x45d6 */
            {8'h00}, /* 0x45d5 */
            {8'h00}, /* 0x45d4 */
            {8'h00}, /* 0x45d3 */
            {8'h00}, /* 0x45d2 */
            {8'h00}, /* 0x45d1 */
            {8'h00}, /* 0x45d0 */
            {8'h00}, /* 0x45cf */
            {8'h00}, /* 0x45ce */
            {8'h00}, /* 0x45cd */
            {8'h00}, /* 0x45cc */
            {8'h00}, /* 0x45cb */
            {8'h00}, /* 0x45ca */
            {8'h00}, /* 0x45c9 */
            {8'h00}, /* 0x45c8 */
            {8'h00}, /* 0x45c7 */
            {8'h00}, /* 0x45c6 */
            {8'h00}, /* 0x45c5 */
            {8'h00}, /* 0x45c4 */
            {8'h00}, /* 0x45c3 */
            {8'h00}, /* 0x45c2 */
            {8'h00}, /* 0x45c1 */
            {8'h00}, /* 0x45c0 */
            {8'h00}, /* 0x45bf */
            {8'h00}, /* 0x45be */
            {8'h00}, /* 0x45bd */
            {8'h00}, /* 0x45bc */
            {8'h00}, /* 0x45bb */
            {8'h00}, /* 0x45ba */
            {8'h00}, /* 0x45b9 */
            {8'h00}, /* 0x45b8 */
            {8'h00}, /* 0x45b7 */
            {8'h00}, /* 0x45b6 */
            {8'h00}, /* 0x45b5 */
            {8'h00}, /* 0x45b4 */
            {8'h00}, /* 0x45b3 */
            {8'h00}, /* 0x45b2 */
            {8'h00}, /* 0x45b1 */
            {8'h00}, /* 0x45b0 */
            {8'h00}, /* 0x45af */
            {8'h00}, /* 0x45ae */
            {8'h00}, /* 0x45ad */
            {8'h00}, /* 0x45ac */
            {8'h00}, /* 0x45ab */
            {8'h00}, /* 0x45aa */
            {8'h00}, /* 0x45a9 */
            {8'h00}, /* 0x45a8 */
            {8'h00}, /* 0x45a7 */
            {8'h00}, /* 0x45a6 */
            {8'h00}, /* 0x45a5 */
            {8'h00}, /* 0x45a4 */
            {8'h00}, /* 0x45a3 */
            {8'h00}, /* 0x45a2 */
            {8'h00}, /* 0x45a1 */
            {8'h00}, /* 0x45a0 */
            {8'h00}, /* 0x459f */
            {8'h00}, /* 0x459e */
            {8'h00}, /* 0x459d */
            {8'h00}, /* 0x459c */
            {8'h00}, /* 0x459b */
            {8'h00}, /* 0x459a */
            {8'h00}, /* 0x4599 */
            {8'h00}, /* 0x4598 */
            {8'h00}, /* 0x4597 */
            {8'h00}, /* 0x4596 */
            {8'h00}, /* 0x4595 */
            {8'h00}, /* 0x4594 */
            {8'h00}, /* 0x4593 */
            {8'h00}, /* 0x4592 */
            {8'h00}, /* 0x4591 */
            {8'h00}, /* 0x4590 */
            {8'h00}, /* 0x458f */
            {8'h00}, /* 0x458e */
            {8'h00}, /* 0x458d */
            {8'h00}, /* 0x458c */
            {8'h00}, /* 0x458b */
            {8'h00}, /* 0x458a */
            {8'h00}, /* 0x4589 */
            {8'h00}, /* 0x4588 */
            {8'h00}, /* 0x4587 */
            {8'h00}, /* 0x4586 */
            {8'h00}, /* 0x4585 */
            {8'h00}, /* 0x4584 */
            {8'h00}, /* 0x4583 */
            {8'h00}, /* 0x4582 */
            {8'h00}, /* 0x4581 */
            {8'h00}, /* 0x4580 */
            {8'h00}, /* 0x457f */
            {8'h00}, /* 0x457e */
            {8'h00}, /* 0x457d */
            {8'h00}, /* 0x457c */
            {8'h00}, /* 0x457b */
            {8'h00}, /* 0x457a */
            {8'h00}, /* 0x4579 */
            {8'h00}, /* 0x4578 */
            {8'h00}, /* 0x4577 */
            {8'h00}, /* 0x4576 */
            {8'h00}, /* 0x4575 */
            {8'h00}, /* 0x4574 */
            {8'h00}, /* 0x4573 */
            {8'h00}, /* 0x4572 */
            {8'h00}, /* 0x4571 */
            {8'h00}, /* 0x4570 */
            {8'h00}, /* 0x456f */
            {8'h00}, /* 0x456e */
            {8'h00}, /* 0x456d */
            {8'h00}, /* 0x456c */
            {8'h00}, /* 0x456b */
            {8'h00}, /* 0x456a */
            {8'h00}, /* 0x4569 */
            {8'h00}, /* 0x4568 */
            {8'h00}, /* 0x4567 */
            {8'h00}, /* 0x4566 */
            {8'h00}, /* 0x4565 */
            {8'h00}, /* 0x4564 */
            {8'h00}, /* 0x4563 */
            {8'h00}, /* 0x4562 */
            {8'h00}, /* 0x4561 */
            {8'h00}, /* 0x4560 */
            {8'h00}, /* 0x455f */
            {8'h00}, /* 0x455e */
            {8'h00}, /* 0x455d */
            {8'h00}, /* 0x455c */
            {8'h00}, /* 0x455b */
            {8'h00}, /* 0x455a */
            {8'h00}, /* 0x4559 */
            {8'h00}, /* 0x4558 */
            {8'h00}, /* 0x4557 */
            {8'h00}, /* 0x4556 */
            {8'h00}, /* 0x4555 */
            {8'h00}, /* 0x4554 */
            {8'h00}, /* 0x4553 */
            {8'h00}, /* 0x4552 */
            {8'h00}, /* 0x4551 */
            {8'h00}, /* 0x4550 */
            {8'h00}, /* 0x454f */
            {8'h00}, /* 0x454e */
            {8'h00}, /* 0x454d */
            {8'h00}, /* 0x454c */
            {8'h00}, /* 0x454b */
            {8'h00}, /* 0x454a */
            {8'h00}, /* 0x4549 */
            {8'h00}, /* 0x4548 */
            {8'h00}, /* 0x4547 */
            {8'h00}, /* 0x4546 */
            {8'h00}, /* 0x4545 */
            {8'h00}, /* 0x4544 */
            {8'h00}, /* 0x4543 */
            {8'h00}, /* 0x4542 */
            {8'h00}, /* 0x4541 */
            {8'h00}, /* 0x4540 */
            {8'h00}, /* 0x453f */
            {8'h00}, /* 0x453e */
            {8'h00}, /* 0x453d */
            {8'h00}, /* 0x453c */
            {8'h00}, /* 0x453b */
            {8'h00}, /* 0x453a */
            {8'h00}, /* 0x4539 */
            {8'h00}, /* 0x4538 */
            {8'h00}, /* 0x4537 */
            {8'h00}, /* 0x4536 */
            {8'h00}, /* 0x4535 */
            {8'h00}, /* 0x4534 */
            {8'h00}, /* 0x4533 */
            {8'h00}, /* 0x4532 */
            {8'h00}, /* 0x4531 */
            {8'h00}, /* 0x4530 */
            {8'h00}, /* 0x452f */
            {8'h00}, /* 0x452e */
            {8'h00}, /* 0x452d */
            {8'h00}, /* 0x452c */
            {8'h00}, /* 0x452b */
            {8'h00}, /* 0x452a */
            {8'h00}, /* 0x4529 */
            {8'h00}, /* 0x4528 */
            {8'h00}, /* 0x4527 */
            {8'h00}, /* 0x4526 */
            {8'h00}, /* 0x4525 */
            {8'h00}, /* 0x4524 */
            {8'h00}, /* 0x4523 */
            {8'h00}, /* 0x4522 */
            {8'h00}, /* 0x4521 */
            {8'h00}, /* 0x4520 */
            {8'h00}, /* 0x451f */
            {8'h00}, /* 0x451e */
            {8'h00}, /* 0x451d */
            {8'h00}, /* 0x451c */
            {8'h00}, /* 0x451b */
            {8'h00}, /* 0x451a */
            {8'h00}, /* 0x4519 */
            {8'h00}, /* 0x4518 */
            {8'h00}, /* 0x4517 */
            {8'h00}, /* 0x4516 */
            {8'h00}, /* 0x4515 */
            {8'h00}, /* 0x4514 */
            {8'h00}, /* 0x4513 */
            {8'h00}, /* 0x4512 */
            {8'h00}, /* 0x4511 */
            {8'h00}, /* 0x4510 */
            {8'h00}, /* 0x450f */
            {8'h00}, /* 0x450e */
            {8'h00}, /* 0x450d */
            {8'h00}, /* 0x450c */
            {8'h00}, /* 0x450b */
            {8'h00}, /* 0x450a */
            {8'h00}, /* 0x4509 */
            {8'h00}, /* 0x4508 */
            {8'h00}, /* 0x4507 */
            {8'h00}, /* 0x4506 */
            {8'h00}, /* 0x4505 */
            {8'h00}, /* 0x4504 */
            {8'h00}, /* 0x4503 */
            {8'h00}, /* 0x4502 */
            {8'h00}, /* 0x4501 */
            {8'h00}, /* 0x4500 */
            {8'h00}, /* 0x44ff */
            {8'h00}, /* 0x44fe */
            {8'h00}, /* 0x44fd */
            {8'h00}, /* 0x44fc */
            {8'h00}, /* 0x44fb */
            {8'h00}, /* 0x44fa */
            {8'h00}, /* 0x44f9 */
            {8'h00}, /* 0x44f8 */
            {8'h00}, /* 0x44f7 */
            {8'h00}, /* 0x44f6 */
            {8'h00}, /* 0x44f5 */
            {8'h00}, /* 0x44f4 */
            {8'h00}, /* 0x44f3 */
            {8'h00}, /* 0x44f2 */
            {8'h00}, /* 0x44f1 */
            {8'h00}, /* 0x44f0 */
            {8'h00}, /* 0x44ef */
            {8'h00}, /* 0x44ee */
            {8'h00}, /* 0x44ed */
            {8'h00}, /* 0x44ec */
            {8'h00}, /* 0x44eb */
            {8'h00}, /* 0x44ea */
            {8'h00}, /* 0x44e9 */
            {8'h00}, /* 0x44e8 */
            {8'h00}, /* 0x44e7 */
            {8'h00}, /* 0x44e6 */
            {8'h00}, /* 0x44e5 */
            {8'h00}, /* 0x44e4 */
            {8'h00}, /* 0x44e3 */
            {8'h00}, /* 0x44e2 */
            {8'h00}, /* 0x44e1 */
            {8'h00}, /* 0x44e0 */
            {8'h00}, /* 0x44df */
            {8'h00}, /* 0x44de */
            {8'h00}, /* 0x44dd */
            {8'h00}, /* 0x44dc */
            {8'h00}, /* 0x44db */
            {8'h00}, /* 0x44da */
            {8'h00}, /* 0x44d9 */
            {8'h00}, /* 0x44d8 */
            {8'h00}, /* 0x44d7 */
            {8'h00}, /* 0x44d6 */
            {8'h00}, /* 0x44d5 */
            {8'h00}, /* 0x44d4 */
            {8'h00}, /* 0x44d3 */
            {8'h00}, /* 0x44d2 */
            {8'h00}, /* 0x44d1 */
            {8'h00}, /* 0x44d0 */
            {8'h00}, /* 0x44cf */
            {8'h00}, /* 0x44ce */
            {8'h00}, /* 0x44cd */
            {8'h00}, /* 0x44cc */
            {8'h00}, /* 0x44cb */
            {8'h00}, /* 0x44ca */
            {8'h00}, /* 0x44c9 */
            {8'h00}, /* 0x44c8 */
            {8'h00}, /* 0x44c7 */
            {8'h00}, /* 0x44c6 */
            {8'h00}, /* 0x44c5 */
            {8'h00}, /* 0x44c4 */
            {8'h00}, /* 0x44c3 */
            {8'h00}, /* 0x44c2 */
            {8'h00}, /* 0x44c1 */
            {8'h00}, /* 0x44c0 */
            {8'h00}, /* 0x44bf */
            {8'h00}, /* 0x44be */
            {8'h00}, /* 0x44bd */
            {8'h00}, /* 0x44bc */
            {8'h00}, /* 0x44bb */
            {8'h00}, /* 0x44ba */
            {8'h00}, /* 0x44b9 */
            {8'h00}, /* 0x44b8 */
            {8'h00}, /* 0x44b7 */
            {8'h00}, /* 0x44b6 */
            {8'h00}, /* 0x44b5 */
            {8'h00}, /* 0x44b4 */
            {8'h00}, /* 0x44b3 */
            {8'h00}, /* 0x44b2 */
            {8'h00}, /* 0x44b1 */
            {8'h00}, /* 0x44b0 */
            {8'h00}, /* 0x44af */
            {8'h00}, /* 0x44ae */
            {8'h00}, /* 0x44ad */
            {8'h00}, /* 0x44ac */
            {8'h00}, /* 0x44ab */
            {8'h00}, /* 0x44aa */
            {8'h00}, /* 0x44a9 */
            {8'h00}, /* 0x44a8 */
            {8'h00}, /* 0x44a7 */
            {8'h00}, /* 0x44a6 */
            {8'h00}, /* 0x44a5 */
            {8'h00}, /* 0x44a4 */
            {8'h00}, /* 0x44a3 */
            {8'h00}, /* 0x44a2 */
            {8'h00}, /* 0x44a1 */
            {8'h00}, /* 0x44a0 */
            {8'h00}, /* 0x449f */
            {8'h00}, /* 0x449e */
            {8'h00}, /* 0x449d */
            {8'h00}, /* 0x449c */
            {8'h00}, /* 0x449b */
            {8'h00}, /* 0x449a */
            {8'h00}, /* 0x4499 */
            {8'h00}, /* 0x4498 */
            {8'h00}, /* 0x4497 */
            {8'h00}, /* 0x4496 */
            {8'h00}, /* 0x4495 */
            {8'h00}, /* 0x4494 */
            {8'h00}, /* 0x4493 */
            {8'h00}, /* 0x4492 */
            {8'h00}, /* 0x4491 */
            {8'h00}, /* 0x4490 */
            {8'h00}, /* 0x448f */
            {8'h00}, /* 0x448e */
            {8'h00}, /* 0x448d */
            {8'h00}, /* 0x448c */
            {8'h00}, /* 0x448b */
            {8'h00}, /* 0x448a */
            {8'h00}, /* 0x4489 */
            {8'h00}, /* 0x4488 */
            {8'h00}, /* 0x4487 */
            {8'h00}, /* 0x4486 */
            {8'h00}, /* 0x4485 */
            {8'h00}, /* 0x4484 */
            {8'h00}, /* 0x4483 */
            {8'h00}, /* 0x4482 */
            {8'h00}, /* 0x4481 */
            {8'h00}, /* 0x4480 */
            {8'h00}, /* 0x447f */
            {8'h00}, /* 0x447e */
            {8'h00}, /* 0x447d */
            {8'h00}, /* 0x447c */
            {8'h00}, /* 0x447b */
            {8'h00}, /* 0x447a */
            {8'h00}, /* 0x4479 */
            {8'h00}, /* 0x4478 */
            {8'h00}, /* 0x4477 */
            {8'h00}, /* 0x4476 */
            {8'h00}, /* 0x4475 */
            {8'h00}, /* 0x4474 */
            {8'h00}, /* 0x4473 */
            {8'h00}, /* 0x4472 */
            {8'h00}, /* 0x4471 */
            {8'h00}, /* 0x4470 */
            {8'h00}, /* 0x446f */
            {8'h00}, /* 0x446e */
            {8'h00}, /* 0x446d */
            {8'h00}, /* 0x446c */
            {8'h00}, /* 0x446b */
            {8'h00}, /* 0x446a */
            {8'h00}, /* 0x4469 */
            {8'h00}, /* 0x4468 */
            {8'h00}, /* 0x4467 */
            {8'h00}, /* 0x4466 */
            {8'h00}, /* 0x4465 */
            {8'h00}, /* 0x4464 */
            {8'h00}, /* 0x4463 */
            {8'h00}, /* 0x4462 */
            {8'h00}, /* 0x4461 */
            {8'h00}, /* 0x4460 */
            {8'h00}, /* 0x445f */
            {8'h00}, /* 0x445e */
            {8'h00}, /* 0x445d */
            {8'h00}, /* 0x445c */
            {8'h00}, /* 0x445b */
            {8'h00}, /* 0x445a */
            {8'h00}, /* 0x4459 */
            {8'h00}, /* 0x4458 */
            {8'h00}, /* 0x4457 */
            {8'h00}, /* 0x4456 */
            {8'h00}, /* 0x4455 */
            {8'h00}, /* 0x4454 */
            {8'h00}, /* 0x4453 */
            {8'h00}, /* 0x4452 */
            {8'h00}, /* 0x4451 */
            {8'h00}, /* 0x4450 */
            {8'h00}, /* 0x444f */
            {8'h00}, /* 0x444e */
            {8'h00}, /* 0x444d */
            {8'h00}, /* 0x444c */
            {8'h00}, /* 0x444b */
            {8'h00}, /* 0x444a */
            {8'h00}, /* 0x4449 */
            {8'h00}, /* 0x4448 */
            {8'h00}, /* 0x4447 */
            {8'h00}, /* 0x4446 */
            {8'h00}, /* 0x4445 */
            {8'h00}, /* 0x4444 */
            {8'h00}, /* 0x4443 */
            {8'h00}, /* 0x4442 */
            {8'h00}, /* 0x4441 */
            {8'h00}, /* 0x4440 */
            {8'h00}, /* 0x443f */
            {8'h00}, /* 0x443e */
            {8'h00}, /* 0x443d */
            {8'h00}, /* 0x443c */
            {8'h00}, /* 0x443b */
            {8'h00}, /* 0x443a */
            {8'h00}, /* 0x4439 */
            {8'h00}, /* 0x4438 */
            {8'h00}, /* 0x4437 */
            {8'h00}, /* 0x4436 */
            {8'h00}, /* 0x4435 */
            {8'h00}, /* 0x4434 */
            {8'h00}, /* 0x4433 */
            {8'h00}, /* 0x4432 */
            {8'h00}, /* 0x4431 */
            {8'h00}, /* 0x4430 */
            {8'h00}, /* 0x442f */
            {8'h00}, /* 0x442e */
            {8'h00}, /* 0x442d */
            {8'h00}, /* 0x442c */
            {8'h00}, /* 0x442b */
            {8'h00}, /* 0x442a */
            {8'h00}, /* 0x4429 */
            {8'h00}, /* 0x4428 */
            {8'h00}, /* 0x4427 */
            {8'h00}, /* 0x4426 */
            {8'h00}, /* 0x4425 */
            {8'h00}, /* 0x4424 */
            {8'h00}, /* 0x4423 */
            {8'h00}, /* 0x4422 */
            {8'h00}, /* 0x4421 */
            {8'h00}, /* 0x4420 */
            {8'h00}, /* 0x441f */
            {8'h00}, /* 0x441e */
            {8'h00}, /* 0x441d */
            {8'h00}, /* 0x441c */
            {8'h00}, /* 0x441b */
            {8'h00}, /* 0x441a */
            {8'h00}, /* 0x4419 */
            {8'h00}, /* 0x4418 */
            {8'h00}, /* 0x4417 */
            {8'h00}, /* 0x4416 */
            {8'h00}, /* 0x4415 */
            {8'h00}, /* 0x4414 */
            {8'h00}, /* 0x4413 */
            {8'h00}, /* 0x4412 */
            {8'h00}, /* 0x4411 */
            {8'h00}, /* 0x4410 */
            {8'h00}, /* 0x440f */
            {8'h00}, /* 0x440e */
            {8'h00}, /* 0x440d */
            {8'h00}, /* 0x440c */
            {8'h00}, /* 0x440b */
            {8'h00}, /* 0x440a */
            {8'h00}, /* 0x4409 */
            {8'h00}, /* 0x4408 */
            {8'h00}, /* 0x4407 */
            {8'h00}, /* 0x4406 */
            {8'h00}, /* 0x4405 */
            {8'h00}, /* 0x4404 */
            {8'h00}, /* 0x4403 */
            {8'h00}, /* 0x4402 */
            {8'h00}, /* 0x4401 */
            {8'h00}, /* 0x4400 */
            {8'h00}, /* 0x43ff */
            {8'h00}, /* 0x43fe */
            {8'h00}, /* 0x43fd */
            {8'h00}, /* 0x43fc */
            {8'h00}, /* 0x43fb */
            {8'h00}, /* 0x43fa */
            {8'h00}, /* 0x43f9 */
            {8'h00}, /* 0x43f8 */
            {8'h00}, /* 0x43f7 */
            {8'h00}, /* 0x43f6 */
            {8'h00}, /* 0x43f5 */
            {8'h00}, /* 0x43f4 */
            {8'h00}, /* 0x43f3 */
            {8'h00}, /* 0x43f2 */
            {8'h00}, /* 0x43f1 */
            {8'h00}, /* 0x43f0 */
            {8'h00}, /* 0x43ef */
            {8'h00}, /* 0x43ee */
            {8'h00}, /* 0x43ed */
            {8'h00}, /* 0x43ec */
            {8'h00}, /* 0x43eb */
            {8'h00}, /* 0x43ea */
            {8'h00}, /* 0x43e9 */
            {8'h00}, /* 0x43e8 */
            {8'h00}, /* 0x43e7 */
            {8'h00}, /* 0x43e6 */
            {8'h00}, /* 0x43e5 */
            {8'h00}, /* 0x43e4 */
            {8'h00}, /* 0x43e3 */
            {8'h00}, /* 0x43e2 */
            {8'h00}, /* 0x43e1 */
            {8'h00}, /* 0x43e0 */
            {8'h00}, /* 0x43df */
            {8'h00}, /* 0x43de */
            {8'h00}, /* 0x43dd */
            {8'h00}, /* 0x43dc */
            {8'h00}, /* 0x43db */
            {8'h00}, /* 0x43da */
            {8'h00}, /* 0x43d9 */
            {8'h00}, /* 0x43d8 */
            {8'h00}, /* 0x43d7 */
            {8'h00}, /* 0x43d6 */
            {8'h00}, /* 0x43d5 */
            {8'h00}, /* 0x43d4 */
            {8'h00}, /* 0x43d3 */
            {8'h00}, /* 0x43d2 */
            {8'h00}, /* 0x43d1 */
            {8'h00}, /* 0x43d0 */
            {8'h00}, /* 0x43cf */
            {8'h00}, /* 0x43ce */
            {8'h00}, /* 0x43cd */
            {8'h00}, /* 0x43cc */
            {8'h00}, /* 0x43cb */
            {8'h00}, /* 0x43ca */
            {8'h00}, /* 0x43c9 */
            {8'h00}, /* 0x43c8 */
            {8'h00}, /* 0x43c7 */
            {8'h00}, /* 0x43c6 */
            {8'h00}, /* 0x43c5 */
            {8'h00}, /* 0x43c4 */
            {8'h00}, /* 0x43c3 */
            {8'h00}, /* 0x43c2 */
            {8'h00}, /* 0x43c1 */
            {8'h00}, /* 0x43c0 */
            {8'h00}, /* 0x43bf */
            {8'h00}, /* 0x43be */
            {8'h00}, /* 0x43bd */
            {8'h00}, /* 0x43bc */
            {8'h00}, /* 0x43bb */
            {8'h00}, /* 0x43ba */
            {8'h00}, /* 0x43b9 */
            {8'h00}, /* 0x43b8 */
            {8'h00}, /* 0x43b7 */
            {8'h00}, /* 0x43b6 */
            {8'h00}, /* 0x43b5 */
            {8'h00}, /* 0x43b4 */
            {8'h00}, /* 0x43b3 */
            {8'h00}, /* 0x43b2 */
            {8'h00}, /* 0x43b1 */
            {8'h00}, /* 0x43b0 */
            {8'h00}, /* 0x43af */
            {8'h00}, /* 0x43ae */
            {8'h00}, /* 0x43ad */
            {8'h00}, /* 0x43ac */
            {8'h00}, /* 0x43ab */
            {8'h00}, /* 0x43aa */
            {8'h00}, /* 0x43a9 */
            {8'h00}, /* 0x43a8 */
            {8'h00}, /* 0x43a7 */
            {8'h00}, /* 0x43a6 */
            {8'h00}, /* 0x43a5 */
            {8'h00}, /* 0x43a4 */
            {8'h00}, /* 0x43a3 */
            {8'h00}, /* 0x43a2 */
            {8'h00}, /* 0x43a1 */
            {8'h00}, /* 0x43a0 */
            {8'h00}, /* 0x439f */
            {8'h00}, /* 0x439e */
            {8'h00}, /* 0x439d */
            {8'h00}, /* 0x439c */
            {8'h00}, /* 0x439b */
            {8'h00}, /* 0x439a */
            {8'h00}, /* 0x4399 */
            {8'h00}, /* 0x4398 */
            {8'h00}, /* 0x4397 */
            {8'h00}, /* 0x4396 */
            {8'h00}, /* 0x4395 */
            {8'h00}, /* 0x4394 */
            {8'h00}, /* 0x4393 */
            {8'h00}, /* 0x4392 */
            {8'h00}, /* 0x4391 */
            {8'h00}, /* 0x4390 */
            {8'h00}, /* 0x438f */
            {8'h00}, /* 0x438e */
            {8'h00}, /* 0x438d */
            {8'h00}, /* 0x438c */
            {8'h00}, /* 0x438b */
            {8'h00}, /* 0x438a */
            {8'h00}, /* 0x4389 */
            {8'h00}, /* 0x4388 */
            {8'h00}, /* 0x4387 */
            {8'h00}, /* 0x4386 */
            {8'h00}, /* 0x4385 */
            {8'h00}, /* 0x4384 */
            {8'h00}, /* 0x4383 */
            {8'h00}, /* 0x4382 */
            {8'h00}, /* 0x4381 */
            {8'h00}, /* 0x4380 */
            {8'h00}, /* 0x437f */
            {8'h00}, /* 0x437e */
            {8'h00}, /* 0x437d */
            {8'h00}, /* 0x437c */
            {8'h00}, /* 0x437b */
            {8'h00}, /* 0x437a */
            {8'h00}, /* 0x4379 */
            {8'h00}, /* 0x4378 */
            {8'h00}, /* 0x4377 */
            {8'h00}, /* 0x4376 */
            {8'h00}, /* 0x4375 */
            {8'h00}, /* 0x4374 */
            {8'h00}, /* 0x4373 */
            {8'h00}, /* 0x4372 */
            {8'h00}, /* 0x4371 */
            {8'h00}, /* 0x4370 */
            {8'h00}, /* 0x436f */
            {8'h00}, /* 0x436e */
            {8'h00}, /* 0x436d */
            {8'h00}, /* 0x436c */
            {8'h00}, /* 0x436b */
            {8'h00}, /* 0x436a */
            {8'h00}, /* 0x4369 */
            {8'h00}, /* 0x4368 */
            {8'h00}, /* 0x4367 */
            {8'h00}, /* 0x4366 */
            {8'h00}, /* 0x4365 */
            {8'h00}, /* 0x4364 */
            {8'h00}, /* 0x4363 */
            {8'h00}, /* 0x4362 */
            {8'h00}, /* 0x4361 */
            {8'h00}, /* 0x4360 */
            {8'h00}, /* 0x435f */
            {8'h00}, /* 0x435e */
            {8'h00}, /* 0x435d */
            {8'h00}, /* 0x435c */
            {8'h00}, /* 0x435b */
            {8'h00}, /* 0x435a */
            {8'h00}, /* 0x4359 */
            {8'h00}, /* 0x4358 */
            {8'h00}, /* 0x4357 */
            {8'h00}, /* 0x4356 */
            {8'h00}, /* 0x4355 */
            {8'h00}, /* 0x4354 */
            {8'h00}, /* 0x4353 */
            {8'h00}, /* 0x4352 */
            {8'h00}, /* 0x4351 */
            {8'h00}, /* 0x4350 */
            {8'h00}, /* 0x434f */
            {8'h00}, /* 0x434e */
            {8'h00}, /* 0x434d */
            {8'h00}, /* 0x434c */
            {8'h00}, /* 0x434b */
            {8'h00}, /* 0x434a */
            {8'h00}, /* 0x4349 */
            {8'h00}, /* 0x4348 */
            {8'h00}, /* 0x4347 */
            {8'h00}, /* 0x4346 */
            {8'h00}, /* 0x4345 */
            {8'h00}, /* 0x4344 */
            {8'h00}, /* 0x4343 */
            {8'h00}, /* 0x4342 */
            {8'h00}, /* 0x4341 */
            {8'h00}, /* 0x4340 */
            {8'h00}, /* 0x433f */
            {8'h00}, /* 0x433e */
            {8'h00}, /* 0x433d */
            {8'h00}, /* 0x433c */
            {8'h00}, /* 0x433b */
            {8'h00}, /* 0x433a */
            {8'h00}, /* 0x4339 */
            {8'h00}, /* 0x4338 */
            {8'h00}, /* 0x4337 */
            {8'h00}, /* 0x4336 */
            {8'h00}, /* 0x4335 */
            {8'h00}, /* 0x4334 */
            {8'h00}, /* 0x4333 */
            {8'h00}, /* 0x4332 */
            {8'h00}, /* 0x4331 */
            {8'h00}, /* 0x4330 */
            {8'h00}, /* 0x432f */
            {8'h00}, /* 0x432e */
            {8'h00}, /* 0x432d */
            {8'h00}, /* 0x432c */
            {8'h00}, /* 0x432b */
            {8'h00}, /* 0x432a */
            {8'h00}, /* 0x4329 */
            {8'h00}, /* 0x4328 */
            {8'h00}, /* 0x4327 */
            {8'h00}, /* 0x4326 */
            {8'h00}, /* 0x4325 */
            {8'h00}, /* 0x4324 */
            {8'h00}, /* 0x4323 */
            {8'h00}, /* 0x4322 */
            {8'h00}, /* 0x4321 */
            {8'h00}, /* 0x4320 */
            {8'h00}, /* 0x431f */
            {8'h00}, /* 0x431e */
            {8'h00}, /* 0x431d */
            {8'h00}, /* 0x431c */
            {8'h00}, /* 0x431b */
            {8'h00}, /* 0x431a */
            {8'h00}, /* 0x4319 */
            {8'h00}, /* 0x4318 */
            {8'h00}, /* 0x4317 */
            {8'h00}, /* 0x4316 */
            {8'h00}, /* 0x4315 */
            {8'h00}, /* 0x4314 */
            {8'h00}, /* 0x4313 */
            {8'h00}, /* 0x4312 */
            {8'h00}, /* 0x4311 */
            {8'h00}, /* 0x4310 */
            {8'h00}, /* 0x430f */
            {8'h00}, /* 0x430e */
            {8'h00}, /* 0x430d */
            {8'h00}, /* 0x430c */
            {8'h00}, /* 0x430b */
            {8'h00}, /* 0x430a */
            {8'h00}, /* 0x4309 */
            {8'h00}, /* 0x4308 */
            {8'h00}, /* 0x4307 */
            {8'h00}, /* 0x4306 */
            {8'h00}, /* 0x4305 */
            {8'h00}, /* 0x4304 */
            {8'h00}, /* 0x4303 */
            {8'h00}, /* 0x4302 */
            {8'h00}, /* 0x4301 */
            {8'h00}, /* 0x4300 */
            {8'h00}, /* 0x42ff */
            {8'h00}, /* 0x42fe */
            {8'h00}, /* 0x42fd */
            {8'h00}, /* 0x42fc */
            {8'h00}, /* 0x42fb */
            {8'h00}, /* 0x42fa */
            {8'h00}, /* 0x42f9 */
            {8'h00}, /* 0x42f8 */
            {8'h00}, /* 0x42f7 */
            {8'h00}, /* 0x42f6 */
            {8'h00}, /* 0x42f5 */
            {8'h00}, /* 0x42f4 */
            {8'h00}, /* 0x42f3 */
            {8'h00}, /* 0x42f2 */
            {8'h00}, /* 0x42f1 */
            {8'h00}, /* 0x42f0 */
            {8'h00}, /* 0x42ef */
            {8'h00}, /* 0x42ee */
            {8'h00}, /* 0x42ed */
            {8'h00}, /* 0x42ec */
            {8'h00}, /* 0x42eb */
            {8'h00}, /* 0x42ea */
            {8'h00}, /* 0x42e9 */
            {8'h00}, /* 0x42e8 */
            {8'h00}, /* 0x42e7 */
            {8'h00}, /* 0x42e6 */
            {8'h00}, /* 0x42e5 */
            {8'h00}, /* 0x42e4 */
            {8'h00}, /* 0x42e3 */
            {8'h00}, /* 0x42e2 */
            {8'h00}, /* 0x42e1 */
            {8'h00}, /* 0x42e0 */
            {8'h00}, /* 0x42df */
            {8'h00}, /* 0x42de */
            {8'h00}, /* 0x42dd */
            {8'h00}, /* 0x42dc */
            {8'h00}, /* 0x42db */
            {8'h00}, /* 0x42da */
            {8'h00}, /* 0x42d9 */
            {8'h00}, /* 0x42d8 */
            {8'h00}, /* 0x42d7 */
            {8'h00}, /* 0x42d6 */
            {8'h00}, /* 0x42d5 */
            {8'h00}, /* 0x42d4 */
            {8'h00}, /* 0x42d3 */
            {8'h00}, /* 0x42d2 */
            {8'h00}, /* 0x42d1 */
            {8'h00}, /* 0x42d0 */
            {8'h00}, /* 0x42cf */
            {8'h00}, /* 0x42ce */
            {8'h00}, /* 0x42cd */
            {8'h00}, /* 0x42cc */
            {8'h00}, /* 0x42cb */
            {8'h00}, /* 0x42ca */
            {8'h00}, /* 0x42c9 */
            {8'h00}, /* 0x42c8 */
            {8'h00}, /* 0x42c7 */
            {8'h00}, /* 0x42c6 */
            {8'h00}, /* 0x42c5 */
            {8'h00}, /* 0x42c4 */
            {8'h00}, /* 0x42c3 */
            {8'h00}, /* 0x42c2 */
            {8'h00}, /* 0x42c1 */
            {8'h00}, /* 0x42c0 */
            {8'h00}, /* 0x42bf */
            {8'h00}, /* 0x42be */
            {8'h00}, /* 0x42bd */
            {8'h00}, /* 0x42bc */
            {8'h00}, /* 0x42bb */
            {8'h00}, /* 0x42ba */
            {8'h00}, /* 0x42b9 */
            {8'h00}, /* 0x42b8 */
            {8'h00}, /* 0x42b7 */
            {8'h00}, /* 0x42b6 */
            {8'h00}, /* 0x42b5 */
            {8'h00}, /* 0x42b4 */
            {8'h00}, /* 0x42b3 */
            {8'h00}, /* 0x42b2 */
            {8'h00}, /* 0x42b1 */
            {8'h00}, /* 0x42b0 */
            {8'h00}, /* 0x42af */
            {8'h00}, /* 0x42ae */
            {8'h00}, /* 0x42ad */
            {8'h00}, /* 0x42ac */
            {8'h00}, /* 0x42ab */
            {8'h00}, /* 0x42aa */
            {8'h00}, /* 0x42a9 */
            {8'h00}, /* 0x42a8 */
            {8'h00}, /* 0x42a7 */
            {8'h00}, /* 0x42a6 */
            {8'h00}, /* 0x42a5 */
            {8'h00}, /* 0x42a4 */
            {8'h00}, /* 0x42a3 */
            {8'h00}, /* 0x42a2 */
            {8'h00}, /* 0x42a1 */
            {8'h00}, /* 0x42a0 */
            {8'h00}, /* 0x429f */
            {8'h00}, /* 0x429e */
            {8'h00}, /* 0x429d */
            {8'h00}, /* 0x429c */
            {8'h00}, /* 0x429b */
            {8'h00}, /* 0x429a */
            {8'h00}, /* 0x4299 */
            {8'h00}, /* 0x4298 */
            {8'h00}, /* 0x4297 */
            {8'h00}, /* 0x4296 */
            {8'h00}, /* 0x4295 */
            {8'h00}, /* 0x4294 */
            {8'h00}, /* 0x4293 */
            {8'h00}, /* 0x4292 */
            {8'h00}, /* 0x4291 */
            {8'h00}, /* 0x4290 */
            {8'h00}, /* 0x428f */
            {8'h00}, /* 0x428e */
            {8'h00}, /* 0x428d */
            {8'h00}, /* 0x428c */
            {8'h00}, /* 0x428b */
            {8'h00}, /* 0x428a */
            {8'h00}, /* 0x4289 */
            {8'h00}, /* 0x4288 */
            {8'h00}, /* 0x4287 */
            {8'h00}, /* 0x4286 */
            {8'h00}, /* 0x4285 */
            {8'h00}, /* 0x4284 */
            {8'h00}, /* 0x4283 */
            {8'h00}, /* 0x4282 */
            {8'h00}, /* 0x4281 */
            {8'h00}, /* 0x4280 */
            {8'h00}, /* 0x427f */
            {8'h00}, /* 0x427e */
            {8'h00}, /* 0x427d */
            {8'h00}, /* 0x427c */
            {8'h00}, /* 0x427b */
            {8'h00}, /* 0x427a */
            {8'h00}, /* 0x4279 */
            {8'h00}, /* 0x4278 */
            {8'h00}, /* 0x4277 */
            {8'h00}, /* 0x4276 */
            {8'h00}, /* 0x4275 */
            {8'h00}, /* 0x4274 */
            {8'h00}, /* 0x4273 */
            {8'h00}, /* 0x4272 */
            {8'h00}, /* 0x4271 */
            {8'h00}, /* 0x4270 */
            {8'h00}, /* 0x426f */
            {8'h00}, /* 0x426e */
            {8'h00}, /* 0x426d */
            {8'h00}, /* 0x426c */
            {8'h00}, /* 0x426b */
            {8'h00}, /* 0x426a */
            {8'h00}, /* 0x4269 */
            {8'h00}, /* 0x4268 */
            {8'h00}, /* 0x4267 */
            {8'h00}, /* 0x4266 */
            {8'h00}, /* 0x4265 */
            {8'h00}, /* 0x4264 */
            {8'h00}, /* 0x4263 */
            {8'h00}, /* 0x4262 */
            {8'h00}, /* 0x4261 */
            {8'h00}, /* 0x4260 */
            {8'h00}, /* 0x425f */
            {8'h00}, /* 0x425e */
            {8'h00}, /* 0x425d */
            {8'h00}, /* 0x425c */
            {8'h00}, /* 0x425b */
            {8'h00}, /* 0x425a */
            {8'h00}, /* 0x4259 */
            {8'h00}, /* 0x4258 */
            {8'h00}, /* 0x4257 */
            {8'h00}, /* 0x4256 */
            {8'h00}, /* 0x4255 */
            {8'h00}, /* 0x4254 */
            {8'h00}, /* 0x4253 */
            {8'h00}, /* 0x4252 */
            {8'h00}, /* 0x4251 */
            {8'h00}, /* 0x4250 */
            {8'h00}, /* 0x424f */
            {8'h00}, /* 0x424e */
            {8'h00}, /* 0x424d */
            {8'h00}, /* 0x424c */
            {8'h00}, /* 0x424b */
            {8'h00}, /* 0x424a */
            {8'h00}, /* 0x4249 */
            {8'h00}, /* 0x4248 */
            {8'h00}, /* 0x4247 */
            {8'h00}, /* 0x4246 */
            {8'h00}, /* 0x4245 */
            {8'h00}, /* 0x4244 */
            {8'h00}, /* 0x4243 */
            {8'h00}, /* 0x4242 */
            {8'h00}, /* 0x4241 */
            {8'h00}, /* 0x4240 */
            {8'h00}, /* 0x423f */
            {8'h00}, /* 0x423e */
            {8'h00}, /* 0x423d */
            {8'h00}, /* 0x423c */
            {8'h00}, /* 0x423b */
            {8'h00}, /* 0x423a */
            {8'h00}, /* 0x4239 */
            {8'h00}, /* 0x4238 */
            {8'h00}, /* 0x4237 */
            {8'h00}, /* 0x4236 */
            {8'h00}, /* 0x4235 */
            {8'h00}, /* 0x4234 */
            {8'h00}, /* 0x4233 */
            {8'h00}, /* 0x4232 */
            {8'h00}, /* 0x4231 */
            {8'h00}, /* 0x4230 */
            {8'h00}, /* 0x422f */
            {8'h00}, /* 0x422e */
            {8'h00}, /* 0x422d */
            {8'h00}, /* 0x422c */
            {8'h00}, /* 0x422b */
            {8'h00}, /* 0x422a */
            {8'h00}, /* 0x4229 */
            {8'h00}, /* 0x4228 */
            {8'h00}, /* 0x4227 */
            {8'h00}, /* 0x4226 */
            {8'h00}, /* 0x4225 */
            {8'h00}, /* 0x4224 */
            {8'h00}, /* 0x4223 */
            {8'h00}, /* 0x4222 */
            {8'h00}, /* 0x4221 */
            {8'h00}, /* 0x4220 */
            {8'h00}, /* 0x421f */
            {8'h00}, /* 0x421e */
            {8'h00}, /* 0x421d */
            {8'h00}, /* 0x421c */
            {8'h00}, /* 0x421b */
            {8'h00}, /* 0x421a */
            {8'h00}, /* 0x4219 */
            {8'h00}, /* 0x4218 */
            {8'h00}, /* 0x4217 */
            {8'h00}, /* 0x4216 */
            {8'h00}, /* 0x4215 */
            {8'h00}, /* 0x4214 */
            {8'h00}, /* 0x4213 */
            {8'h00}, /* 0x4212 */
            {8'h00}, /* 0x4211 */
            {8'h00}, /* 0x4210 */
            {8'h00}, /* 0x420f */
            {8'h00}, /* 0x420e */
            {8'h00}, /* 0x420d */
            {8'h00}, /* 0x420c */
            {8'h00}, /* 0x420b */
            {8'h00}, /* 0x420a */
            {8'h00}, /* 0x4209 */
            {8'h00}, /* 0x4208 */
            {8'h00}, /* 0x4207 */
            {8'h00}, /* 0x4206 */
            {8'h00}, /* 0x4205 */
            {8'h00}, /* 0x4204 */
            {8'h00}, /* 0x4203 */
            {8'h00}, /* 0x4202 */
            {8'h00}, /* 0x4201 */
            {8'h00}, /* 0x4200 */
            {8'h00}, /* 0x41ff */
            {8'h00}, /* 0x41fe */
            {8'h00}, /* 0x41fd */
            {8'h00}, /* 0x41fc */
            {8'h00}, /* 0x41fb */
            {8'h00}, /* 0x41fa */
            {8'h00}, /* 0x41f9 */
            {8'h00}, /* 0x41f8 */
            {8'h00}, /* 0x41f7 */
            {8'h00}, /* 0x41f6 */
            {8'h00}, /* 0x41f5 */
            {8'h00}, /* 0x41f4 */
            {8'h00}, /* 0x41f3 */
            {8'h00}, /* 0x41f2 */
            {8'h00}, /* 0x41f1 */
            {8'h00}, /* 0x41f0 */
            {8'h00}, /* 0x41ef */
            {8'h00}, /* 0x41ee */
            {8'h00}, /* 0x41ed */
            {8'h00}, /* 0x41ec */
            {8'h00}, /* 0x41eb */
            {8'h00}, /* 0x41ea */
            {8'h00}, /* 0x41e9 */
            {8'h00}, /* 0x41e8 */
            {8'h00}, /* 0x41e7 */
            {8'h00}, /* 0x41e6 */
            {8'h00}, /* 0x41e5 */
            {8'h00}, /* 0x41e4 */
            {8'h00}, /* 0x41e3 */
            {8'h00}, /* 0x41e2 */
            {8'h00}, /* 0x41e1 */
            {8'h00}, /* 0x41e0 */
            {8'h00}, /* 0x41df */
            {8'h00}, /* 0x41de */
            {8'h00}, /* 0x41dd */
            {8'h00}, /* 0x41dc */
            {8'h00}, /* 0x41db */
            {8'h00}, /* 0x41da */
            {8'h00}, /* 0x41d9 */
            {8'h00}, /* 0x41d8 */
            {8'h00}, /* 0x41d7 */
            {8'h00}, /* 0x41d6 */
            {8'h00}, /* 0x41d5 */
            {8'h00}, /* 0x41d4 */
            {8'h00}, /* 0x41d3 */
            {8'h00}, /* 0x41d2 */
            {8'h00}, /* 0x41d1 */
            {8'h00}, /* 0x41d0 */
            {8'h00}, /* 0x41cf */
            {8'h00}, /* 0x41ce */
            {8'h00}, /* 0x41cd */
            {8'h00}, /* 0x41cc */
            {8'h00}, /* 0x41cb */
            {8'h00}, /* 0x41ca */
            {8'h00}, /* 0x41c9 */
            {8'h00}, /* 0x41c8 */
            {8'h00}, /* 0x41c7 */
            {8'h00}, /* 0x41c6 */
            {8'h00}, /* 0x41c5 */
            {8'h00}, /* 0x41c4 */
            {8'h00}, /* 0x41c3 */
            {8'h00}, /* 0x41c2 */
            {8'h00}, /* 0x41c1 */
            {8'h00}, /* 0x41c0 */
            {8'h00}, /* 0x41bf */
            {8'h00}, /* 0x41be */
            {8'h00}, /* 0x41bd */
            {8'h00}, /* 0x41bc */
            {8'h00}, /* 0x41bb */
            {8'h00}, /* 0x41ba */
            {8'h00}, /* 0x41b9 */
            {8'h00}, /* 0x41b8 */
            {8'h00}, /* 0x41b7 */
            {8'h00}, /* 0x41b6 */
            {8'h00}, /* 0x41b5 */
            {8'h00}, /* 0x41b4 */
            {8'h00}, /* 0x41b3 */
            {8'h00}, /* 0x41b2 */
            {8'h00}, /* 0x41b1 */
            {8'h00}, /* 0x41b0 */
            {8'h00}, /* 0x41af */
            {8'h00}, /* 0x41ae */
            {8'h00}, /* 0x41ad */
            {8'h00}, /* 0x41ac */
            {8'h00}, /* 0x41ab */
            {8'h00}, /* 0x41aa */
            {8'h00}, /* 0x41a9 */
            {8'h00}, /* 0x41a8 */
            {8'h00}, /* 0x41a7 */
            {8'h00}, /* 0x41a6 */
            {8'h00}, /* 0x41a5 */
            {8'h00}, /* 0x41a4 */
            {8'h00}, /* 0x41a3 */
            {8'h00}, /* 0x41a2 */
            {8'h00}, /* 0x41a1 */
            {8'h00}, /* 0x41a0 */
            {8'h00}, /* 0x419f */
            {8'h00}, /* 0x419e */
            {8'h00}, /* 0x419d */
            {8'h00}, /* 0x419c */
            {8'h00}, /* 0x419b */
            {8'h00}, /* 0x419a */
            {8'h00}, /* 0x4199 */
            {8'h00}, /* 0x4198 */
            {8'h00}, /* 0x4197 */
            {8'h00}, /* 0x4196 */
            {8'h00}, /* 0x4195 */
            {8'h00}, /* 0x4194 */
            {8'h00}, /* 0x4193 */
            {8'h00}, /* 0x4192 */
            {8'h00}, /* 0x4191 */
            {8'h00}, /* 0x4190 */
            {8'h00}, /* 0x418f */
            {8'h00}, /* 0x418e */
            {8'h00}, /* 0x418d */
            {8'h00}, /* 0x418c */
            {8'h00}, /* 0x418b */
            {8'h00}, /* 0x418a */
            {8'h00}, /* 0x4189 */
            {8'h00}, /* 0x4188 */
            {8'h00}, /* 0x4187 */
            {8'h00}, /* 0x4186 */
            {8'h00}, /* 0x4185 */
            {8'h00}, /* 0x4184 */
            {8'h00}, /* 0x4183 */
            {8'h00}, /* 0x4182 */
            {8'h00}, /* 0x4181 */
            {8'h00}, /* 0x4180 */
            {8'h00}, /* 0x417f */
            {8'h00}, /* 0x417e */
            {8'h00}, /* 0x417d */
            {8'h00}, /* 0x417c */
            {8'h00}, /* 0x417b */
            {8'h00}, /* 0x417a */
            {8'h00}, /* 0x4179 */
            {8'h00}, /* 0x4178 */
            {8'h00}, /* 0x4177 */
            {8'h00}, /* 0x4176 */
            {8'h00}, /* 0x4175 */
            {8'h00}, /* 0x4174 */
            {8'h00}, /* 0x4173 */
            {8'h00}, /* 0x4172 */
            {8'h00}, /* 0x4171 */
            {8'h00}, /* 0x4170 */
            {8'h00}, /* 0x416f */
            {8'h00}, /* 0x416e */
            {8'h00}, /* 0x416d */
            {8'h00}, /* 0x416c */
            {8'h00}, /* 0x416b */
            {8'h00}, /* 0x416a */
            {8'h00}, /* 0x4169 */
            {8'h00}, /* 0x4168 */
            {8'h00}, /* 0x4167 */
            {8'h00}, /* 0x4166 */
            {8'h00}, /* 0x4165 */
            {8'h00}, /* 0x4164 */
            {8'h00}, /* 0x4163 */
            {8'h00}, /* 0x4162 */
            {8'h00}, /* 0x4161 */
            {8'h00}, /* 0x4160 */
            {8'h00}, /* 0x415f */
            {8'h00}, /* 0x415e */
            {8'h00}, /* 0x415d */
            {8'h00}, /* 0x415c */
            {8'h00}, /* 0x415b */
            {8'h00}, /* 0x415a */
            {8'h00}, /* 0x4159 */
            {8'h00}, /* 0x4158 */
            {8'h00}, /* 0x4157 */
            {8'h00}, /* 0x4156 */
            {8'h00}, /* 0x4155 */
            {8'h00}, /* 0x4154 */
            {8'h00}, /* 0x4153 */
            {8'h00}, /* 0x4152 */
            {8'h00}, /* 0x4151 */
            {8'h00}, /* 0x4150 */
            {8'h00}, /* 0x414f */
            {8'h00}, /* 0x414e */
            {8'h00}, /* 0x414d */
            {8'h00}, /* 0x414c */
            {8'h00}, /* 0x414b */
            {8'h00}, /* 0x414a */
            {8'h00}, /* 0x4149 */
            {8'h00}, /* 0x4148 */
            {8'h00}, /* 0x4147 */
            {8'h00}, /* 0x4146 */
            {8'h00}, /* 0x4145 */
            {8'h00}, /* 0x4144 */
            {8'h00}, /* 0x4143 */
            {8'h00}, /* 0x4142 */
            {8'h00}, /* 0x4141 */
            {8'h00}, /* 0x4140 */
            {8'h00}, /* 0x413f */
            {8'h00}, /* 0x413e */
            {8'h00}, /* 0x413d */
            {8'h00}, /* 0x413c */
            {8'h00}, /* 0x413b */
            {8'h00}, /* 0x413a */
            {8'h00}, /* 0x4139 */
            {8'h00}, /* 0x4138 */
            {8'h00}, /* 0x4137 */
            {8'h00}, /* 0x4136 */
            {8'h00}, /* 0x4135 */
            {8'h00}, /* 0x4134 */
            {8'h00}, /* 0x4133 */
            {8'h00}, /* 0x4132 */
            {8'h00}, /* 0x4131 */
            {8'h00}, /* 0x4130 */
            {8'h00}, /* 0x412f */
            {8'h00}, /* 0x412e */
            {8'h00}, /* 0x412d */
            {8'h00}, /* 0x412c */
            {8'h00}, /* 0x412b */
            {8'h00}, /* 0x412a */
            {8'h00}, /* 0x4129 */
            {8'h00}, /* 0x4128 */
            {8'h00}, /* 0x4127 */
            {8'h00}, /* 0x4126 */
            {8'h00}, /* 0x4125 */
            {8'h00}, /* 0x4124 */
            {8'h00}, /* 0x4123 */
            {8'h00}, /* 0x4122 */
            {8'h00}, /* 0x4121 */
            {8'h00}, /* 0x4120 */
            {8'h00}, /* 0x411f */
            {8'h00}, /* 0x411e */
            {8'h00}, /* 0x411d */
            {8'h00}, /* 0x411c */
            {8'h00}, /* 0x411b */
            {8'h00}, /* 0x411a */
            {8'h00}, /* 0x4119 */
            {8'h00}, /* 0x4118 */
            {8'h00}, /* 0x4117 */
            {8'h00}, /* 0x4116 */
            {8'h00}, /* 0x4115 */
            {8'h00}, /* 0x4114 */
            {8'h00}, /* 0x4113 */
            {8'h00}, /* 0x4112 */
            {8'h00}, /* 0x4111 */
            {8'h00}, /* 0x4110 */
            {8'h00}, /* 0x410f */
            {8'h00}, /* 0x410e */
            {8'h00}, /* 0x410d */
            {8'h00}, /* 0x410c */
            {8'h00}, /* 0x410b */
            {8'h00}, /* 0x410a */
            {8'h00}, /* 0x4109 */
            {8'h00}, /* 0x4108 */
            {8'h00}, /* 0x4107 */
            {8'h00}, /* 0x4106 */
            {8'h00}, /* 0x4105 */
            {8'h00}, /* 0x4104 */
            {8'h00}, /* 0x4103 */
            {8'h00}, /* 0x4102 */
            {8'h00}, /* 0x4101 */
            {8'h00}, /* 0x4100 */
            {8'h00}, /* 0x40ff */
            {8'h00}, /* 0x40fe */
            {8'h00}, /* 0x40fd */
            {8'h00}, /* 0x40fc */
            {8'h00}, /* 0x40fb */
            {8'h00}, /* 0x40fa */
            {8'h00}, /* 0x40f9 */
            {8'h00}, /* 0x40f8 */
            {8'h00}, /* 0x40f7 */
            {8'h00}, /* 0x40f6 */
            {8'h00}, /* 0x40f5 */
            {8'h00}, /* 0x40f4 */
            {8'h00}, /* 0x40f3 */
            {8'h00}, /* 0x40f2 */
            {8'h00}, /* 0x40f1 */
            {8'h00}, /* 0x40f0 */
            {8'h00}, /* 0x40ef */
            {8'h00}, /* 0x40ee */
            {8'h00}, /* 0x40ed */
            {8'h00}, /* 0x40ec */
            {8'h00}, /* 0x40eb */
            {8'h00}, /* 0x40ea */
            {8'h00}, /* 0x40e9 */
            {8'h00}, /* 0x40e8 */
            {8'h00}, /* 0x40e7 */
            {8'h00}, /* 0x40e6 */
            {8'h00}, /* 0x40e5 */
            {8'h00}, /* 0x40e4 */
            {8'h00}, /* 0x40e3 */
            {8'h00}, /* 0x40e2 */
            {8'h00}, /* 0x40e1 */
            {8'h00}, /* 0x40e0 */
            {8'h00}, /* 0x40df */
            {8'h00}, /* 0x40de */
            {8'h00}, /* 0x40dd */
            {8'h00}, /* 0x40dc */
            {8'h00}, /* 0x40db */
            {8'h00}, /* 0x40da */
            {8'h00}, /* 0x40d9 */
            {8'h00}, /* 0x40d8 */
            {8'h00}, /* 0x40d7 */
            {8'h00}, /* 0x40d6 */
            {8'h00}, /* 0x40d5 */
            {8'h00}, /* 0x40d4 */
            {8'h00}, /* 0x40d3 */
            {8'h00}, /* 0x40d2 */
            {8'h00}, /* 0x40d1 */
            {8'h00}, /* 0x40d0 */
            {8'h00}, /* 0x40cf */
            {8'h00}, /* 0x40ce */
            {8'h00}, /* 0x40cd */
            {8'h00}, /* 0x40cc */
            {8'h00}, /* 0x40cb */
            {8'h00}, /* 0x40ca */
            {8'h00}, /* 0x40c9 */
            {8'h00}, /* 0x40c8 */
            {8'h00}, /* 0x40c7 */
            {8'h00}, /* 0x40c6 */
            {8'h00}, /* 0x40c5 */
            {8'h00}, /* 0x40c4 */
            {8'h00}, /* 0x40c3 */
            {8'h00}, /* 0x40c2 */
            {8'h00}, /* 0x40c1 */
            {8'h00}, /* 0x40c0 */
            {8'h00}, /* 0x40bf */
            {8'h00}, /* 0x40be */
            {8'h00}, /* 0x40bd */
            {8'h00}, /* 0x40bc */
            {8'h00}, /* 0x40bb */
            {8'h00}, /* 0x40ba */
            {8'h00}, /* 0x40b9 */
            {8'h00}, /* 0x40b8 */
            {8'h00}, /* 0x40b7 */
            {8'h00}, /* 0x40b6 */
            {8'h00}, /* 0x40b5 */
            {8'h00}, /* 0x40b4 */
            {8'h00}, /* 0x40b3 */
            {8'h00}, /* 0x40b2 */
            {8'h00}, /* 0x40b1 */
            {8'h00}, /* 0x40b0 */
            {8'h00}, /* 0x40af */
            {8'h00}, /* 0x40ae */
            {8'h00}, /* 0x40ad */
            {8'h00}, /* 0x40ac */
            {8'h00}, /* 0x40ab */
            {8'h00}, /* 0x40aa */
            {8'h00}, /* 0x40a9 */
            {8'h00}, /* 0x40a8 */
            {8'h00}, /* 0x40a7 */
            {8'h00}, /* 0x40a6 */
            {8'h00}, /* 0x40a5 */
            {8'h00}, /* 0x40a4 */
            {8'h00}, /* 0x40a3 */
            {8'h00}, /* 0x40a2 */
            {8'h00}, /* 0x40a1 */
            {8'h00}, /* 0x40a0 */
            {8'h00}, /* 0x409f */
            {8'h00}, /* 0x409e */
            {8'h00}, /* 0x409d */
            {8'h00}, /* 0x409c */
            {8'h00}, /* 0x409b */
            {8'h00}, /* 0x409a */
            {8'h00}, /* 0x4099 */
            {8'h00}, /* 0x4098 */
            {8'h00}, /* 0x4097 */
            {8'h00}, /* 0x4096 */
            {8'h00}, /* 0x4095 */
            {8'h00}, /* 0x4094 */
            {8'h00}, /* 0x4093 */
            {8'h00}, /* 0x4092 */
            {8'h00}, /* 0x4091 */
            {8'h00}, /* 0x4090 */
            {8'h00}, /* 0x408f */
            {8'h00}, /* 0x408e */
            {8'h00}, /* 0x408d */
            {8'h00}, /* 0x408c */
            {8'h00}, /* 0x408b */
            {8'h00}, /* 0x408a */
            {8'h00}, /* 0x4089 */
            {8'h00}, /* 0x4088 */
            {8'h00}, /* 0x4087 */
            {8'h00}, /* 0x4086 */
            {8'h00}, /* 0x4085 */
            {8'h00}, /* 0x4084 */
            {8'h00}, /* 0x4083 */
            {8'h00}, /* 0x4082 */
            {8'h00}, /* 0x4081 */
            {8'h00}, /* 0x4080 */
            {8'h00}, /* 0x407f */
            {8'h00}, /* 0x407e */
            {8'h00}, /* 0x407d */
            {8'h00}, /* 0x407c */
            {8'h00}, /* 0x407b */
            {8'h00}, /* 0x407a */
            {8'h00}, /* 0x4079 */
            {8'h00}, /* 0x4078 */
            {8'h00}, /* 0x4077 */
            {8'h00}, /* 0x4076 */
            {8'h00}, /* 0x4075 */
            {8'h00}, /* 0x4074 */
            {8'h00}, /* 0x4073 */
            {8'h00}, /* 0x4072 */
            {8'h00}, /* 0x4071 */
            {8'h00}, /* 0x4070 */
            {8'h00}, /* 0x406f */
            {8'h00}, /* 0x406e */
            {8'h00}, /* 0x406d */
            {8'h00}, /* 0x406c */
            {8'h00}, /* 0x406b */
            {8'h00}, /* 0x406a */
            {8'h00}, /* 0x4069 */
            {8'h00}, /* 0x4068 */
            {8'h00}, /* 0x4067 */
            {8'h00}, /* 0x4066 */
            {8'h00}, /* 0x4065 */
            {8'h00}, /* 0x4064 */
            {8'h00}, /* 0x4063 */
            {8'h00}, /* 0x4062 */
            {8'h00}, /* 0x4061 */
            {8'h00}, /* 0x4060 */
            {8'h00}, /* 0x405f */
            {8'h00}, /* 0x405e */
            {8'h00}, /* 0x405d */
            {8'h00}, /* 0x405c */
            {8'h00}, /* 0x405b */
            {8'h00}, /* 0x405a */
            {8'h00}, /* 0x4059 */
            {8'h00}, /* 0x4058 */
            {8'h00}, /* 0x4057 */
            {8'h00}, /* 0x4056 */
            {8'h00}, /* 0x4055 */
            {8'h00}, /* 0x4054 */
            {8'h00}, /* 0x4053 */
            {8'h00}, /* 0x4052 */
            {8'h00}, /* 0x4051 */
            {8'h00}, /* 0x4050 */
            {8'h00}, /* 0x404f */
            {8'h00}, /* 0x404e */
            {8'h00}, /* 0x404d */
            {8'h00}, /* 0x404c */
            {8'h00}, /* 0x404b */
            {8'h00}, /* 0x404a */
            {8'h00}, /* 0x4049 */
            {8'h00}, /* 0x4048 */
            {8'h00}, /* 0x4047 */
            {8'h00}, /* 0x4046 */
            {8'h00}, /* 0x4045 */
            {8'h00}, /* 0x4044 */
            {8'h00}, /* 0x4043 */
            {8'h00}, /* 0x4042 */
            {8'h00}, /* 0x4041 */
            {8'h00}, /* 0x4040 */
            {8'h00}, /* 0x403f */
            {8'h00}, /* 0x403e */
            {8'h00}, /* 0x403d */
            {8'h00}, /* 0x403c */
            {8'h00}, /* 0x403b */
            {8'h00}, /* 0x403a */
            {8'h00}, /* 0x4039 */
            {8'h00}, /* 0x4038 */
            {8'h00}, /* 0x4037 */
            {8'h00}, /* 0x4036 */
            {8'h00}, /* 0x4035 */
            {8'h00}, /* 0x4034 */
            {8'h00}, /* 0x4033 */
            {8'h00}, /* 0x4032 */
            {8'h00}, /* 0x4031 */
            {8'h00}, /* 0x4030 */
            {8'h00}, /* 0x402f */
            {8'h00}, /* 0x402e */
            {8'h00}, /* 0x402d */
            {8'h00}, /* 0x402c */
            {8'h00}, /* 0x402b */
            {8'h00}, /* 0x402a */
            {8'h00}, /* 0x4029 */
            {8'h00}, /* 0x4028 */
            {8'h00}, /* 0x4027 */
            {8'h00}, /* 0x4026 */
            {8'h00}, /* 0x4025 */
            {8'h00}, /* 0x4024 */
            {8'h00}, /* 0x4023 */
            {8'h00}, /* 0x4022 */
            {8'h00}, /* 0x4021 */
            {8'h00}, /* 0x4020 */
            {8'h00}, /* 0x401f */
            {8'h00}, /* 0x401e */
            {8'h00}, /* 0x401d */
            {8'h00}, /* 0x401c */
            {8'h00}, /* 0x401b */
            {8'h00}, /* 0x401a */
            {8'h00}, /* 0x4019 */
            {8'h00}, /* 0x4018 */
            {8'h00}, /* 0x4017 */
            {8'h00}, /* 0x4016 */
            {8'h00}, /* 0x4015 */
            {8'h00}, /* 0x4014 */
            {8'h00}, /* 0x4013 */
            {8'h00}, /* 0x4012 */
            {8'h00}, /* 0x4011 */
            {8'h00}, /* 0x4010 */
            {8'h00}, /* 0x400f */
            {8'h00}, /* 0x400e */
            {8'h00}, /* 0x400d */
            {8'h00}, /* 0x400c */
            {8'h00}, /* 0x400b */
            {8'h00}, /* 0x400a */
            {8'h00}, /* 0x4009 */
            {8'h00}, /* 0x4008 */
            {8'h00}, /* 0x4007 */
            {8'h00}, /* 0x4006 */
            {8'h00}, /* 0x4005 */
            {8'h00}, /* 0x4004 */
            {8'h00}, /* 0x4003 */
            {8'h00}, /* 0x4002 */
            {8'h00}, /* 0x4001 */
            {8'h00}, /* 0x4000 */
            {8'h00}, /* 0x3fff */
            {8'h00}, /* 0x3ffe */
            {8'h00}, /* 0x3ffd */
            {8'h00}, /* 0x3ffc */
            {8'h00}, /* 0x3ffb */
            {8'h00}, /* 0x3ffa */
            {8'h00}, /* 0x3ff9 */
            {8'h00}, /* 0x3ff8 */
            {8'h00}, /* 0x3ff7 */
            {8'h00}, /* 0x3ff6 */
            {8'h00}, /* 0x3ff5 */
            {8'h00}, /* 0x3ff4 */
            {8'h00}, /* 0x3ff3 */
            {8'h00}, /* 0x3ff2 */
            {8'h00}, /* 0x3ff1 */
            {8'h00}, /* 0x3ff0 */
            {8'h00}, /* 0x3fef */
            {8'h00}, /* 0x3fee */
            {8'h00}, /* 0x3fed */
            {8'h00}, /* 0x3fec */
            {8'h00}, /* 0x3feb */
            {8'h00}, /* 0x3fea */
            {8'h00}, /* 0x3fe9 */
            {8'h00}, /* 0x3fe8 */
            {8'h00}, /* 0x3fe7 */
            {8'h00}, /* 0x3fe6 */
            {8'h00}, /* 0x3fe5 */
            {8'h00}, /* 0x3fe4 */
            {8'h00}, /* 0x3fe3 */
            {8'h00}, /* 0x3fe2 */
            {8'h00}, /* 0x3fe1 */
            {8'h00}, /* 0x3fe0 */
            {8'h00}, /* 0x3fdf */
            {8'h00}, /* 0x3fde */
            {8'h00}, /* 0x3fdd */
            {8'h00}, /* 0x3fdc */
            {8'h00}, /* 0x3fdb */
            {8'h00}, /* 0x3fda */
            {8'h00}, /* 0x3fd9 */
            {8'h00}, /* 0x3fd8 */
            {8'h00}, /* 0x3fd7 */
            {8'h00}, /* 0x3fd6 */
            {8'h00}, /* 0x3fd5 */
            {8'h00}, /* 0x3fd4 */
            {8'h00}, /* 0x3fd3 */
            {8'h00}, /* 0x3fd2 */
            {8'h00}, /* 0x3fd1 */
            {8'h00}, /* 0x3fd0 */
            {8'h00}, /* 0x3fcf */
            {8'h00}, /* 0x3fce */
            {8'h00}, /* 0x3fcd */
            {8'h00}, /* 0x3fcc */
            {8'h00}, /* 0x3fcb */
            {8'h00}, /* 0x3fca */
            {8'h00}, /* 0x3fc9 */
            {8'h00}, /* 0x3fc8 */
            {8'h00}, /* 0x3fc7 */
            {8'h00}, /* 0x3fc6 */
            {8'h00}, /* 0x3fc5 */
            {8'h00}, /* 0x3fc4 */
            {8'h00}, /* 0x3fc3 */
            {8'h00}, /* 0x3fc2 */
            {8'h00}, /* 0x3fc1 */
            {8'h00}, /* 0x3fc0 */
            {8'h00}, /* 0x3fbf */
            {8'h00}, /* 0x3fbe */
            {8'h00}, /* 0x3fbd */
            {8'h00}, /* 0x3fbc */
            {8'h00}, /* 0x3fbb */
            {8'h00}, /* 0x3fba */
            {8'h00}, /* 0x3fb9 */
            {8'h00}, /* 0x3fb8 */
            {8'h00}, /* 0x3fb7 */
            {8'h00}, /* 0x3fb6 */
            {8'h00}, /* 0x3fb5 */
            {8'h00}, /* 0x3fb4 */
            {8'h00}, /* 0x3fb3 */
            {8'h00}, /* 0x3fb2 */
            {8'h00}, /* 0x3fb1 */
            {8'h00}, /* 0x3fb0 */
            {8'h00}, /* 0x3faf */
            {8'h00}, /* 0x3fae */
            {8'h00}, /* 0x3fad */
            {8'h00}, /* 0x3fac */
            {8'h00}, /* 0x3fab */
            {8'h00}, /* 0x3faa */
            {8'h00}, /* 0x3fa9 */
            {8'h00}, /* 0x3fa8 */
            {8'h00}, /* 0x3fa7 */
            {8'h00}, /* 0x3fa6 */
            {8'h00}, /* 0x3fa5 */
            {8'h00}, /* 0x3fa4 */
            {8'h00}, /* 0x3fa3 */
            {8'h00}, /* 0x3fa2 */
            {8'h00}, /* 0x3fa1 */
            {8'h00}, /* 0x3fa0 */
            {8'h00}, /* 0x3f9f */
            {8'h00}, /* 0x3f9e */
            {8'h00}, /* 0x3f9d */
            {8'h00}, /* 0x3f9c */
            {8'h00}, /* 0x3f9b */
            {8'h00}, /* 0x3f9a */
            {8'h00}, /* 0x3f99 */
            {8'h00}, /* 0x3f98 */
            {8'h00}, /* 0x3f97 */
            {8'h00}, /* 0x3f96 */
            {8'h00}, /* 0x3f95 */
            {8'h00}, /* 0x3f94 */
            {8'h00}, /* 0x3f93 */
            {8'h00}, /* 0x3f92 */
            {8'h00}, /* 0x3f91 */
            {8'h00}, /* 0x3f90 */
            {8'h00}, /* 0x3f8f */
            {8'h00}, /* 0x3f8e */
            {8'h00}, /* 0x3f8d */
            {8'h00}, /* 0x3f8c */
            {8'h00}, /* 0x3f8b */
            {8'h00}, /* 0x3f8a */
            {8'h00}, /* 0x3f89 */
            {8'h00}, /* 0x3f88 */
            {8'h00}, /* 0x3f87 */
            {8'h00}, /* 0x3f86 */
            {8'h00}, /* 0x3f85 */
            {8'h00}, /* 0x3f84 */
            {8'h00}, /* 0x3f83 */
            {8'h00}, /* 0x3f82 */
            {8'h00}, /* 0x3f81 */
            {8'h00}, /* 0x3f80 */
            {8'h00}, /* 0x3f7f */
            {8'h00}, /* 0x3f7e */
            {8'h00}, /* 0x3f7d */
            {8'h00}, /* 0x3f7c */
            {8'h00}, /* 0x3f7b */
            {8'h00}, /* 0x3f7a */
            {8'h00}, /* 0x3f79 */
            {8'h00}, /* 0x3f78 */
            {8'h00}, /* 0x3f77 */
            {8'h00}, /* 0x3f76 */
            {8'h00}, /* 0x3f75 */
            {8'h00}, /* 0x3f74 */
            {8'h00}, /* 0x3f73 */
            {8'h00}, /* 0x3f72 */
            {8'h00}, /* 0x3f71 */
            {8'h00}, /* 0x3f70 */
            {8'h00}, /* 0x3f6f */
            {8'h00}, /* 0x3f6e */
            {8'h00}, /* 0x3f6d */
            {8'h00}, /* 0x3f6c */
            {8'h00}, /* 0x3f6b */
            {8'h00}, /* 0x3f6a */
            {8'h00}, /* 0x3f69 */
            {8'h00}, /* 0x3f68 */
            {8'h00}, /* 0x3f67 */
            {8'h00}, /* 0x3f66 */
            {8'h00}, /* 0x3f65 */
            {8'h00}, /* 0x3f64 */
            {8'h00}, /* 0x3f63 */
            {8'h00}, /* 0x3f62 */
            {8'h00}, /* 0x3f61 */
            {8'h00}, /* 0x3f60 */
            {8'h00}, /* 0x3f5f */
            {8'h00}, /* 0x3f5e */
            {8'h00}, /* 0x3f5d */
            {8'h00}, /* 0x3f5c */
            {8'h00}, /* 0x3f5b */
            {8'h00}, /* 0x3f5a */
            {8'h00}, /* 0x3f59 */
            {8'h00}, /* 0x3f58 */
            {8'h00}, /* 0x3f57 */
            {8'h00}, /* 0x3f56 */
            {8'h00}, /* 0x3f55 */
            {8'h00}, /* 0x3f54 */
            {8'h00}, /* 0x3f53 */
            {8'h00}, /* 0x3f52 */
            {8'h00}, /* 0x3f51 */
            {8'h00}, /* 0x3f50 */
            {8'h00}, /* 0x3f4f */
            {8'h00}, /* 0x3f4e */
            {8'h00}, /* 0x3f4d */
            {8'h00}, /* 0x3f4c */
            {8'h00}, /* 0x3f4b */
            {8'h00}, /* 0x3f4a */
            {8'h00}, /* 0x3f49 */
            {8'h00}, /* 0x3f48 */
            {8'h00}, /* 0x3f47 */
            {8'h00}, /* 0x3f46 */
            {8'h00}, /* 0x3f45 */
            {8'h00}, /* 0x3f44 */
            {8'h00}, /* 0x3f43 */
            {8'h00}, /* 0x3f42 */
            {8'h00}, /* 0x3f41 */
            {8'h00}, /* 0x3f40 */
            {8'h00}, /* 0x3f3f */
            {8'h00}, /* 0x3f3e */
            {8'h00}, /* 0x3f3d */
            {8'h00}, /* 0x3f3c */
            {8'h00}, /* 0x3f3b */
            {8'h00}, /* 0x3f3a */
            {8'h00}, /* 0x3f39 */
            {8'h00}, /* 0x3f38 */
            {8'h00}, /* 0x3f37 */
            {8'h00}, /* 0x3f36 */
            {8'h00}, /* 0x3f35 */
            {8'h00}, /* 0x3f34 */
            {8'h00}, /* 0x3f33 */
            {8'h00}, /* 0x3f32 */
            {8'h00}, /* 0x3f31 */
            {8'h00}, /* 0x3f30 */
            {8'h00}, /* 0x3f2f */
            {8'h00}, /* 0x3f2e */
            {8'h00}, /* 0x3f2d */
            {8'h00}, /* 0x3f2c */
            {8'h00}, /* 0x3f2b */
            {8'h00}, /* 0x3f2a */
            {8'h00}, /* 0x3f29 */
            {8'h00}, /* 0x3f28 */
            {8'h00}, /* 0x3f27 */
            {8'h00}, /* 0x3f26 */
            {8'h00}, /* 0x3f25 */
            {8'h00}, /* 0x3f24 */
            {8'h00}, /* 0x3f23 */
            {8'h00}, /* 0x3f22 */
            {8'h00}, /* 0x3f21 */
            {8'h00}, /* 0x3f20 */
            {8'h00}, /* 0x3f1f */
            {8'h00}, /* 0x3f1e */
            {8'h00}, /* 0x3f1d */
            {8'h00}, /* 0x3f1c */
            {8'h00}, /* 0x3f1b */
            {8'h00}, /* 0x3f1a */
            {8'h00}, /* 0x3f19 */
            {8'h00}, /* 0x3f18 */
            {8'h00}, /* 0x3f17 */
            {8'h00}, /* 0x3f16 */
            {8'h00}, /* 0x3f15 */
            {8'h00}, /* 0x3f14 */
            {8'h00}, /* 0x3f13 */
            {8'h00}, /* 0x3f12 */
            {8'h00}, /* 0x3f11 */
            {8'h00}, /* 0x3f10 */
            {8'h00}, /* 0x3f0f */
            {8'h00}, /* 0x3f0e */
            {8'h00}, /* 0x3f0d */
            {8'h00}, /* 0x3f0c */
            {8'h00}, /* 0x3f0b */
            {8'h00}, /* 0x3f0a */
            {8'h00}, /* 0x3f09 */
            {8'h00}, /* 0x3f08 */
            {8'h00}, /* 0x3f07 */
            {8'h00}, /* 0x3f06 */
            {8'h00}, /* 0x3f05 */
            {8'h00}, /* 0x3f04 */
            {8'h00}, /* 0x3f03 */
            {8'h00}, /* 0x3f02 */
            {8'h00}, /* 0x3f01 */
            {8'h00}, /* 0x3f00 */
            {8'h00}, /* 0x3eff */
            {8'h00}, /* 0x3efe */
            {8'h00}, /* 0x3efd */
            {8'h00}, /* 0x3efc */
            {8'h00}, /* 0x3efb */
            {8'h00}, /* 0x3efa */
            {8'h00}, /* 0x3ef9 */
            {8'h00}, /* 0x3ef8 */
            {8'h00}, /* 0x3ef7 */
            {8'h00}, /* 0x3ef6 */
            {8'h00}, /* 0x3ef5 */
            {8'h00}, /* 0x3ef4 */
            {8'h00}, /* 0x3ef3 */
            {8'h00}, /* 0x3ef2 */
            {8'h00}, /* 0x3ef1 */
            {8'h00}, /* 0x3ef0 */
            {8'h00}, /* 0x3eef */
            {8'h00}, /* 0x3eee */
            {8'h00}, /* 0x3eed */
            {8'h00}, /* 0x3eec */
            {8'h00}, /* 0x3eeb */
            {8'h00}, /* 0x3eea */
            {8'h00}, /* 0x3ee9 */
            {8'h00}, /* 0x3ee8 */
            {8'h00}, /* 0x3ee7 */
            {8'h00}, /* 0x3ee6 */
            {8'h00}, /* 0x3ee5 */
            {8'h00}, /* 0x3ee4 */
            {8'h00}, /* 0x3ee3 */
            {8'h00}, /* 0x3ee2 */
            {8'h00}, /* 0x3ee1 */
            {8'h00}, /* 0x3ee0 */
            {8'h00}, /* 0x3edf */
            {8'h00}, /* 0x3ede */
            {8'h00}, /* 0x3edd */
            {8'h00}, /* 0x3edc */
            {8'h00}, /* 0x3edb */
            {8'h00}, /* 0x3eda */
            {8'h00}, /* 0x3ed9 */
            {8'h00}, /* 0x3ed8 */
            {8'h00}, /* 0x3ed7 */
            {8'h00}, /* 0x3ed6 */
            {8'h00}, /* 0x3ed5 */
            {8'h00}, /* 0x3ed4 */
            {8'h00}, /* 0x3ed3 */
            {8'h00}, /* 0x3ed2 */
            {8'h00}, /* 0x3ed1 */
            {8'h00}, /* 0x3ed0 */
            {8'h00}, /* 0x3ecf */
            {8'h00}, /* 0x3ece */
            {8'h00}, /* 0x3ecd */
            {8'h00}, /* 0x3ecc */
            {8'h00}, /* 0x3ecb */
            {8'h00}, /* 0x3eca */
            {8'h00}, /* 0x3ec9 */
            {8'h00}, /* 0x3ec8 */
            {8'h00}, /* 0x3ec7 */
            {8'h00}, /* 0x3ec6 */
            {8'h00}, /* 0x3ec5 */
            {8'h00}, /* 0x3ec4 */
            {8'h00}, /* 0x3ec3 */
            {8'h00}, /* 0x3ec2 */
            {8'h00}, /* 0x3ec1 */
            {8'h00}, /* 0x3ec0 */
            {8'h00}, /* 0x3ebf */
            {8'h00}, /* 0x3ebe */
            {8'h00}, /* 0x3ebd */
            {8'h00}, /* 0x3ebc */
            {8'h00}, /* 0x3ebb */
            {8'h00}, /* 0x3eba */
            {8'h00}, /* 0x3eb9 */
            {8'h00}, /* 0x3eb8 */
            {8'h00}, /* 0x3eb7 */
            {8'h00}, /* 0x3eb6 */
            {8'h00}, /* 0x3eb5 */
            {8'h00}, /* 0x3eb4 */
            {8'h00}, /* 0x3eb3 */
            {8'h00}, /* 0x3eb2 */
            {8'h00}, /* 0x3eb1 */
            {8'h00}, /* 0x3eb0 */
            {8'h00}, /* 0x3eaf */
            {8'h00}, /* 0x3eae */
            {8'h00}, /* 0x3ead */
            {8'h00}, /* 0x3eac */
            {8'h00}, /* 0x3eab */
            {8'h00}, /* 0x3eaa */
            {8'h00}, /* 0x3ea9 */
            {8'h00}, /* 0x3ea8 */
            {8'h00}, /* 0x3ea7 */
            {8'h00}, /* 0x3ea6 */
            {8'h00}, /* 0x3ea5 */
            {8'h00}, /* 0x3ea4 */
            {8'h00}, /* 0x3ea3 */
            {8'h00}, /* 0x3ea2 */
            {8'h00}, /* 0x3ea1 */
            {8'h00}, /* 0x3ea0 */
            {8'h00}, /* 0x3e9f */
            {8'h00}, /* 0x3e9e */
            {8'h00}, /* 0x3e9d */
            {8'h00}, /* 0x3e9c */
            {8'h00}, /* 0x3e9b */
            {8'h00}, /* 0x3e9a */
            {8'h00}, /* 0x3e99 */
            {8'h00}, /* 0x3e98 */
            {8'h00}, /* 0x3e97 */
            {8'h00}, /* 0x3e96 */
            {8'h00}, /* 0x3e95 */
            {8'h00}, /* 0x3e94 */
            {8'h00}, /* 0x3e93 */
            {8'h00}, /* 0x3e92 */
            {8'h00}, /* 0x3e91 */
            {8'h00}, /* 0x3e90 */
            {8'h00}, /* 0x3e8f */
            {8'h00}, /* 0x3e8e */
            {8'h00}, /* 0x3e8d */
            {8'h00}, /* 0x3e8c */
            {8'h00}, /* 0x3e8b */
            {8'h00}, /* 0x3e8a */
            {8'h00}, /* 0x3e89 */
            {8'h00}, /* 0x3e88 */
            {8'h00}, /* 0x3e87 */
            {8'h00}, /* 0x3e86 */
            {8'h00}, /* 0x3e85 */
            {8'h00}, /* 0x3e84 */
            {8'h00}, /* 0x3e83 */
            {8'h00}, /* 0x3e82 */
            {8'h00}, /* 0x3e81 */
            {8'h00}, /* 0x3e80 */
            {8'h00}, /* 0x3e7f */
            {8'h00}, /* 0x3e7e */
            {8'h00}, /* 0x3e7d */
            {8'h00}, /* 0x3e7c */
            {8'h00}, /* 0x3e7b */
            {8'h00}, /* 0x3e7a */
            {8'h00}, /* 0x3e79 */
            {8'h00}, /* 0x3e78 */
            {8'h00}, /* 0x3e77 */
            {8'h00}, /* 0x3e76 */
            {8'h00}, /* 0x3e75 */
            {8'h00}, /* 0x3e74 */
            {8'h00}, /* 0x3e73 */
            {8'h00}, /* 0x3e72 */
            {8'h00}, /* 0x3e71 */
            {8'h00}, /* 0x3e70 */
            {8'h00}, /* 0x3e6f */
            {8'h00}, /* 0x3e6e */
            {8'h00}, /* 0x3e6d */
            {8'h00}, /* 0x3e6c */
            {8'h00}, /* 0x3e6b */
            {8'h00}, /* 0x3e6a */
            {8'h00}, /* 0x3e69 */
            {8'h00}, /* 0x3e68 */
            {8'h00}, /* 0x3e67 */
            {8'h00}, /* 0x3e66 */
            {8'h00}, /* 0x3e65 */
            {8'h00}, /* 0x3e64 */
            {8'h00}, /* 0x3e63 */
            {8'h00}, /* 0x3e62 */
            {8'h00}, /* 0x3e61 */
            {8'h00}, /* 0x3e60 */
            {8'h00}, /* 0x3e5f */
            {8'h00}, /* 0x3e5e */
            {8'h00}, /* 0x3e5d */
            {8'h00}, /* 0x3e5c */
            {8'h00}, /* 0x3e5b */
            {8'h00}, /* 0x3e5a */
            {8'h00}, /* 0x3e59 */
            {8'h00}, /* 0x3e58 */
            {8'h00}, /* 0x3e57 */
            {8'h00}, /* 0x3e56 */
            {8'h00}, /* 0x3e55 */
            {8'h00}, /* 0x3e54 */
            {8'h00}, /* 0x3e53 */
            {8'h00}, /* 0x3e52 */
            {8'h00}, /* 0x3e51 */
            {8'h00}, /* 0x3e50 */
            {8'h00}, /* 0x3e4f */
            {8'h00}, /* 0x3e4e */
            {8'h00}, /* 0x3e4d */
            {8'h00}, /* 0x3e4c */
            {8'h00}, /* 0x3e4b */
            {8'h00}, /* 0x3e4a */
            {8'h00}, /* 0x3e49 */
            {8'h00}, /* 0x3e48 */
            {8'h00}, /* 0x3e47 */
            {8'h00}, /* 0x3e46 */
            {8'h00}, /* 0x3e45 */
            {8'h00}, /* 0x3e44 */
            {8'h00}, /* 0x3e43 */
            {8'h00}, /* 0x3e42 */
            {8'h00}, /* 0x3e41 */
            {8'h00}, /* 0x3e40 */
            {8'h00}, /* 0x3e3f */
            {8'h00}, /* 0x3e3e */
            {8'h00}, /* 0x3e3d */
            {8'h00}, /* 0x3e3c */
            {8'h00}, /* 0x3e3b */
            {8'h00}, /* 0x3e3a */
            {8'h00}, /* 0x3e39 */
            {8'h00}, /* 0x3e38 */
            {8'h00}, /* 0x3e37 */
            {8'h00}, /* 0x3e36 */
            {8'h00}, /* 0x3e35 */
            {8'h00}, /* 0x3e34 */
            {8'h00}, /* 0x3e33 */
            {8'h00}, /* 0x3e32 */
            {8'h00}, /* 0x3e31 */
            {8'h00}, /* 0x3e30 */
            {8'h00}, /* 0x3e2f */
            {8'h00}, /* 0x3e2e */
            {8'h00}, /* 0x3e2d */
            {8'h00}, /* 0x3e2c */
            {8'h00}, /* 0x3e2b */
            {8'h00}, /* 0x3e2a */
            {8'h00}, /* 0x3e29 */
            {8'h00}, /* 0x3e28 */
            {8'h00}, /* 0x3e27 */
            {8'h00}, /* 0x3e26 */
            {8'h00}, /* 0x3e25 */
            {8'h00}, /* 0x3e24 */
            {8'h00}, /* 0x3e23 */
            {8'h00}, /* 0x3e22 */
            {8'h00}, /* 0x3e21 */
            {8'h00}, /* 0x3e20 */
            {8'h00}, /* 0x3e1f */
            {8'h00}, /* 0x3e1e */
            {8'h00}, /* 0x3e1d */
            {8'h00}, /* 0x3e1c */
            {8'h00}, /* 0x3e1b */
            {8'h00}, /* 0x3e1a */
            {8'h00}, /* 0x3e19 */
            {8'h00}, /* 0x3e18 */
            {8'h00}, /* 0x3e17 */
            {8'h00}, /* 0x3e16 */
            {8'h00}, /* 0x3e15 */
            {8'h00}, /* 0x3e14 */
            {8'h00}, /* 0x3e13 */
            {8'h00}, /* 0x3e12 */
            {8'h00}, /* 0x3e11 */
            {8'h00}, /* 0x3e10 */
            {8'h00}, /* 0x3e0f */
            {8'h00}, /* 0x3e0e */
            {8'h00}, /* 0x3e0d */
            {8'h00}, /* 0x3e0c */
            {8'h00}, /* 0x3e0b */
            {8'h00}, /* 0x3e0a */
            {8'h00}, /* 0x3e09 */
            {8'h00}, /* 0x3e08 */
            {8'h00}, /* 0x3e07 */
            {8'h00}, /* 0x3e06 */
            {8'h00}, /* 0x3e05 */
            {8'h00}, /* 0x3e04 */
            {8'h00}, /* 0x3e03 */
            {8'h00}, /* 0x3e02 */
            {8'h00}, /* 0x3e01 */
            {8'h00}, /* 0x3e00 */
            {8'h00}, /* 0x3dff */
            {8'h00}, /* 0x3dfe */
            {8'h00}, /* 0x3dfd */
            {8'h00}, /* 0x3dfc */
            {8'h00}, /* 0x3dfb */
            {8'h00}, /* 0x3dfa */
            {8'h00}, /* 0x3df9 */
            {8'h00}, /* 0x3df8 */
            {8'h00}, /* 0x3df7 */
            {8'h00}, /* 0x3df6 */
            {8'h00}, /* 0x3df5 */
            {8'h00}, /* 0x3df4 */
            {8'h00}, /* 0x3df3 */
            {8'h00}, /* 0x3df2 */
            {8'h00}, /* 0x3df1 */
            {8'h00}, /* 0x3df0 */
            {8'h00}, /* 0x3def */
            {8'h00}, /* 0x3dee */
            {8'h00}, /* 0x3ded */
            {8'h00}, /* 0x3dec */
            {8'h00}, /* 0x3deb */
            {8'h00}, /* 0x3dea */
            {8'h00}, /* 0x3de9 */
            {8'h00}, /* 0x3de8 */
            {8'h00}, /* 0x3de7 */
            {8'h00}, /* 0x3de6 */
            {8'h00}, /* 0x3de5 */
            {8'h00}, /* 0x3de4 */
            {8'h00}, /* 0x3de3 */
            {8'h00}, /* 0x3de2 */
            {8'h00}, /* 0x3de1 */
            {8'h00}, /* 0x3de0 */
            {8'h00}, /* 0x3ddf */
            {8'h00}, /* 0x3dde */
            {8'h00}, /* 0x3ddd */
            {8'h00}, /* 0x3ddc */
            {8'h00}, /* 0x3ddb */
            {8'h00}, /* 0x3dda */
            {8'h00}, /* 0x3dd9 */
            {8'h00}, /* 0x3dd8 */
            {8'h00}, /* 0x3dd7 */
            {8'h00}, /* 0x3dd6 */
            {8'h00}, /* 0x3dd5 */
            {8'h00}, /* 0x3dd4 */
            {8'h00}, /* 0x3dd3 */
            {8'h00}, /* 0x3dd2 */
            {8'h00}, /* 0x3dd1 */
            {8'h00}, /* 0x3dd0 */
            {8'h00}, /* 0x3dcf */
            {8'h00}, /* 0x3dce */
            {8'h00}, /* 0x3dcd */
            {8'h00}, /* 0x3dcc */
            {8'h00}, /* 0x3dcb */
            {8'h00}, /* 0x3dca */
            {8'h00}, /* 0x3dc9 */
            {8'h00}, /* 0x3dc8 */
            {8'h00}, /* 0x3dc7 */
            {8'h00}, /* 0x3dc6 */
            {8'h00}, /* 0x3dc5 */
            {8'h00}, /* 0x3dc4 */
            {8'h00}, /* 0x3dc3 */
            {8'h00}, /* 0x3dc2 */
            {8'h00}, /* 0x3dc1 */
            {8'h00}, /* 0x3dc0 */
            {8'h00}, /* 0x3dbf */
            {8'h00}, /* 0x3dbe */
            {8'h00}, /* 0x3dbd */
            {8'h00}, /* 0x3dbc */
            {8'h00}, /* 0x3dbb */
            {8'h00}, /* 0x3dba */
            {8'h00}, /* 0x3db9 */
            {8'h00}, /* 0x3db8 */
            {8'h00}, /* 0x3db7 */
            {8'h00}, /* 0x3db6 */
            {8'h00}, /* 0x3db5 */
            {8'h00}, /* 0x3db4 */
            {8'h00}, /* 0x3db3 */
            {8'h00}, /* 0x3db2 */
            {8'h00}, /* 0x3db1 */
            {8'h00}, /* 0x3db0 */
            {8'h00}, /* 0x3daf */
            {8'h00}, /* 0x3dae */
            {8'h00}, /* 0x3dad */
            {8'h00}, /* 0x3dac */
            {8'h00}, /* 0x3dab */
            {8'h00}, /* 0x3daa */
            {8'h00}, /* 0x3da9 */
            {8'h00}, /* 0x3da8 */
            {8'h00}, /* 0x3da7 */
            {8'h00}, /* 0x3da6 */
            {8'h00}, /* 0x3da5 */
            {8'h00}, /* 0x3da4 */
            {8'h00}, /* 0x3da3 */
            {8'h00}, /* 0x3da2 */
            {8'h00}, /* 0x3da1 */
            {8'h00}, /* 0x3da0 */
            {8'h00}, /* 0x3d9f */
            {8'h00}, /* 0x3d9e */
            {8'h00}, /* 0x3d9d */
            {8'h00}, /* 0x3d9c */
            {8'h00}, /* 0x3d9b */
            {8'h00}, /* 0x3d9a */
            {8'h00}, /* 0x3d99 */
            {8'h00}, /* 0x3d98 */
            {8'h00}, /* 0x3d97 */
            {8'h00}, /* 0x3d96 */
            {8'h00}, /* 0x3d95 */
            {8'h00}, /* 0x3d94 */
            {8'h00}, /* 0x3d93 */
            {8'h00}, /* 0x3d92 */
            {8'h00}, /* 0x3d91 */
            {8'h00}, /* 0x3d90 */
            {8'h00}, /* 0x3d8f */
            {8'h00}, /* 0x3d8e */
            {8'h00}, /* 0x3d8d */
            {8'h00}, /* 0x3d8c */
            {8'h00}, /* 0x3d8b */
            {8'h00}, /* 0x3d8a */
            {8'h00}, /* 0x3d89 */
            {8'h00}, /* 0x3d88 */
            {8'h00}, /* 0x3d87 */
            {8'h00}, /* 0x3d86 */
            {8'h00}, /* 0x3d85 */
            {8'h00}, /* 0x3d84 */
            {8'h00}, /* 0x3d83 */
            {8'h00}, /* 0x3d82 */
            {8'h00}, /* 0x3d81 */
            {8'h00}, /* 0x3d80 */
            {8'h00}, /* 0x3d7f */
            {8'h00}, /* 0x3d7e */
            {8'h00}, /* 0x3d7d */
            {8'h00}, /* 0x3d7c */
            {8'h00}, /* 0x3d7b */
            {8'h00}, /* 0x3d7a */
            {8'h00}, /* 0x3d79 */
            {8'h00}, /* 0x3d78 */
            {8'h00}, /* 0x3d77 */
            {8'h00}, /* 0x3d76 */
            {8'h00}, /* 0x3d75 */
            {8'h00}, /* 0x3d74 */
            {8'h00}, /* 0x3d73 */
            {8'h00}, /* 0x3d72 */
            {8'h00}, /* 0x3d71 */
            {8'h00}, /* 0x3d70 */
            {8'h00}, /* 0x3d6f */
            {8'h00}, /* 0x3d6e */
            {8'h00}, /* 0x3d6d */
            {8'h00}, /* 0x3d6c */
            {8'h00}, /* 0x3d6b */
            {8'h00}, /* 0x3d6a */
            {8'h00}, /* 0x3d69 */
            {8'h00}, /* 0x3d68 */
            {8'h00}, /* 0x3d67 */
            {8'h00}, /* 0x3d66 */
            {8'h00}, /* 0x3d65 */
            {8'h00}, /* 0x3d64 */
            {8'h00}, /* 0x3d63 */
            {8'h00}, /* 0x3d62 */
            {8'h00}, /* 0x3d61 */
            {8'h00}, /* 0x3d60 */
            {8'h00}, /* 0x3d5f */
            {8'h00}, /* 0x3d5e */
            {8'h00}, /* 0x3d5d */
            {8'h00}, /* 0x3d5c */
            {8'h00}, /* 0x3d5b */
            {8'h00}, /* 0x3d5a */
            {8'h00}, /* 0x3d59 */
            {8'h00}, /* 0x3d58 */
            {8'h00}, /* 0x3d57 */
            {8'h00}, /* 0x3d56 */
            {8'h00}, /* 0x3d55 */
            {8'h00}, /* 0x3d54 */
            {8'h00}, /* 0x3d53 */
            {8'h00}, /* 0x3d52 */
            {8'h00}, /* 0x3d51 */
            {8'h00}, /* 0x3d50 */
            {8'h00}, /* 0x3d4f */
            {8'h00}, /* 0x3d4e */
            {8'h00}, /* 0x3d4d */
            {8'h00}, /* 0x3d4c */
            {8'h00}, /* 0x3d4b */
            {8'h00}, /* 0x3d4a */
            {8'h00}, /* 0x3d49 */
            {8'h00}, /* 0x3d48 */
            {8'h00}, /* 0x3d47 */
            {8'h00}, /* 0x3d46 */
            {8'h00}, /* 0x3d45 */
            {8'h00}, /* 0x3d44 */
            {8'h00}, /* 0x3d43 */
            {8'h00}, /* 0x3d42 */
            {8'h00}, /* 0x3d41 */
            {8'h00}, /* 0x3d40 */
            {8'h00}, /* 0x3d3f */
            {8'h00}, /* 0x3d3e */
            {8'h00}, /* 0x3d3d */
            {8'h00}, /* 0x3d3c */
            {8'h00}, /* 0x3d3b */
            {8'h00}, /* 0x3d3a */
            {8'h00}, /* 0x3d39 */
            {8'h00}, /* 0x3d38 */
            {8'h00}, /* 0x3d37 */
            {8'h00}, /* 0x3d36 */
            {8'h00}, /* 0x3d35 */
            {8'h00}, /* 0x3d34 */
            {8'h00}, /* 0x3d33 */
            {8'h00}, /* 0x3d32 */
            {8'h00}, /* 0x3d31 */
            {8'h00}, /* 0x3d30 */
            {8'h00}, /* 0x3d2f */
            {8'h00}, /* 0x3d2e */
            {8'h00}, /* 0x3d2d */
            {8'h00}, /* 0x3d2c */
            {8'h00}, /* 0x3d2b */
            {8'h00}, /* 0x3d2a */
            {8'h00}, /* 0x3d29 */
            {8'h00}, /* 0x3d28 */
            {8'h00}, /* 0x3d27 */
            {8'h00}, /* 0x3d26 */
            {8'h00}, /* 0x3d25 */
            {8'h00}, /* 0x3d24 */
            {8'h00}, /* 0x3d23 */
            {8'h00}, /* 0x3d22 */
            {8'h00}, /* 0x3d21 */
            {8'h00}, /* 0x3d20 */
            {8'h00}, /* 0x3d1f */
            {8'h00}, /* 0x3d1e */
            {8'h00}, /* 0x3d1d */
            {8'h00}, /* 0x3d1c */
            {8'h00}, /* 0x3d1b */
            {8'h00}, /* 0x3d1a */
            {8'h00}, /* 0x3d19 */
            {8'h00}, /* 0x3d18 */
            {8'h00}, /* 0x3d17 */
            {8'h00}, /* 0x3d16 */
            {8'h00}, /* 0x3d15 */
            {8'h00}, /* 0x3d14 */
            {8'h00}, /* 0x3d13 */
            {8'h00}, /* 0x3d12 */
            {8'h00}, /* 0x3d11 */
            {8'h00}, /* 0x3d10 */
            {8'h00}, /* 0x3d0f */
            {8'h00}, /* 0x3d0e */
            {8'h00}, /* 0x3d0d */
            {8'h00}, /* 0x3d0c */
            {8'h00}, /* 0x3d0b */
            {8'h00}, /* 0x3d0a */
            {8'h00}, /* 0x3d09 */
            {8'h00}, /* 0x3d08 */
            {8'h00}, /* 0x3d07 */
            {8'h00}, /* 0x3d06 */
            {8'h00}, /* 0x3d05 */
            {8'h00}, /* 0x3d04 */
            {8'h00}, /* 0x3d03 */
            {8'h00}, /* 0x3d02 */
            {8'h00}, /* 0x3d01 */
            {8'h00}, /* 0x3d00 */
            {8'h00}, /* 0x3cff */
            {8'h00}, /* 0x3cfe */
            {8'h00}, /* 0x3cfd */
            {8'h00}, /* 0x3cfc */
            {8'h00}, /* 0x3cfb */
            {8'h00}, /* 0x3cfa */
            {8'h00}, /* 0x3cf9 */
            {8'h00}, /* 0x3cf8 */
            {8'h00}, /* 0x3cf7 */
            {8'h00}, /* 0x3cf6 */
            {8'h00}, /* 0x3cf5 */
            {8'h00}, /* 0x3cf4 */
            {8'h00}, /* 0x3cf3 */
            {8'h00}, /* 0x3cf2 */
            {8'h00}, /* 0x3cf1 */
            {8'h00}, /* 0x3cf0 */
            {8'h00}, /* 0x3cef */
            {8'h00}, /* 0x3cee */
            {8'h00}, /* 0x3ced */
            {8'h00}, /* 0x3cec */
            {8'h00}, /* 0x3ceb */
            {8'h00}, /* 0x3cea */
            {8'h00}, /* 0x3ce9 */
            {8'h00}, /* 0x3ce8 */
            {8'h00}, /* 0x3ce7 */
            {8'h00}, /* 0x3ce6 */
            {8'h00}, /* 0x3ce5 */
            {8'h00}, /* 0x3ce4 */
            {8'h00}, /* 0x3ce3 */
            {8'h00}, /* 0x3ce2 */
            {8'h00}, /* 0x3ce1 */
            {8'h00}, /* 0x3ce0 */
            {8'h00}, /* 0x3cdf */
            {8'h00}, /* 0x3cde */
            {8'h00}, /* 0x3cdd */
            {8'h00}, /* 0x3cdc */
            {8'h00}, /* 0x3cdb */
            {8'h00}, /* 0x3cda */
            {8'h00}, /* 0x3cd9 */
            {8'h00}, /* 0x3cd8 */
            {8'h00}, /* 0x3cd7 */
            {8'h00}, /* 0x3cd6 */
            {8'h00}, /* 0x3cd5 */
            {8'h00}, /* 0x3cd4 */
            {8'h00}, /* 0x3cd3 */
            {8'h00}, /* 0x3cd2 */
            {8'h00}, /* 0x3cd1 */
            {8'h00}, /* 0x3cd0 */
            {8'h00}, /* 0x3ccf */
            {8'h00}, /* 0x3cce */
            {8'h00}, /* 0x3ccd */
            {8'h00}, /* 0x3ccc */
            {8'h00}, /* 0x3ccb */
            {8'h00}, /* 0x3cca */
            {8'h00}, /* 0x3cc9 */
            {8'h00}, /* 0x3cc8 */
            {8'h00}, /* 0x3cc7 */
            {8'h00}, /* 0x3cc6 */
            {8'h00}, /* 0x3cc5 */
            {8'h00}, /* 0x3cc4 */
            {8'h00}, /* 0x3cc3 */
            {8'h00}, /* 0x3cc2 */
            {8'h00}, /* 0x3cc1 */
            {8'h00}, /* 0x3cc0 */
            {8'h00}, /* 0x3cbf */
            {8'h00}, /* 0x3cbe */
            {8'h00}, /* 0x3cbd */
            {8'h00}, /* 0x3cbc */
            {8'h00}, /* 0x3cbb */
            {8'h00}, /* 0x3cba */
            {8'h00}, /* 0x3cb9 */
            {8'h00}, /* 0x3cb8 */
            {8'h00}, /* 0x3cb7 */
            {8'h00}, /* 0x3cb6 */
            {8'h00}, /* 0x3cb5 */
            {8'h00}, /* 0x3cb4 */
            {8'h00}, /* 0x3cb3 */
            {8'h00}, /* 0x3cb2 */
            {8'h00}, /* 0x3cb1 */
            {8'h00}, /* 0x3cb0 */
            {8'h00}, /* 0x3caf */
            {8'h00}, /* 0x3cae */
            {8'h00}, /* 0x3cad */
            {8'h00}, /* 0x3cac */
            {8'h00}, /* 0x3cab */
            {8'h00}, /* 0x3caa */
            {8'h00}, /* 0x3ca9 */
            {8'h00}, /* 0x3ca8 */
            {8'h00}, /* 0x3ca7 */
            {8'h00}, /* 0x3ca6 */
            {8'h00}, /* 0x3ca5 */
            {8'h00}, /* 0x3ca4 */
            {8'h00}, /* 0x3ca3 */
            {8'h00}, /* 0x3ca2 */
            {8'h00}, /* 0x3ca1 */
            {8'h00}, /* 0x3ca0 */
            {8'h00}, /* 0x3c9f */
            {8'h00}, /* 0x3c9e */
            {8'h00}, /* 0x3c9d */
            {8'h00}, /* 0x3c9c */
            {8'h00}, /* 0x3c9b */
            {8'h00}, /* 0x3c9a */
            {8'h00}, /* 0x3c99 */
            {8'h00}, /* 0x3c98 */
            {8'h00}, /* 0x3c97 */
            {8'h00}, /* 0x3c96 */
            {8'h00}, /* 0x3c95 */
            {8'h00}, /* 0x3c94 */
            {8'h00}, /* 0x3c93 */
            {8'h00}, /* 0x3c92 */
            {8'h00}, /* 0x3c91 */
            {8'h00}, /* 0x3c90 */
            {8'h00}, /* 0x3c8f */
            {8'h00}, /* 0x3c8e */
            {8'h00}, /* 0x3c8d */
            {8'h00}, /* 0x3c8c */
            {8'h00}, /* 0x3c8b */
            {8'h00}, /* 0x3c8a */
            {8'h00}, /* 0x3c89 */
            {8'h00}, /* 0x3c88 */
            {8'h00}, /* 0x3c87 */
            {8'h00}, /* 0x3c86 */
            {8'h00}, /* 0x3c85 */
            {8'h00}, /* 0x3c84 */
            {8'h00}, /* 0x3c83 */
            {8'h00}, /* 0x3c82 */
            {8'h00}, /* 0x3c81 */
            {8'h00}, /* 0x3c80 */
            {8'h00}, /* 0x3c7f */
            {8'h00}, /* 0x3c7e */
            {8'h00}, /* 0x3c7d */
            {8'h00}, /* 0x3c7c */
            {8'h00}, /* 0x3c7b */
            {8'h00}, /* 0x3c7a */
            {8'h00}, /* 0x3c79 */
            {8'h00}, /* 0x3c78 */
            {8'h00}, /* 0x3c77 */
            {8'h00}, /* 0x3c76 */
            {8'h00}, /* 0x3c75 */
            {8'h00}, /* 0x3c74 */
            {8'h00}, /* 0x3c73 */
            {8'h00}, /* 0x3c72 */
            {8'h00}, /* 0x3c71 */
            {8'h00}, /* 0x3c70 */
            {8'h00}, /* 0x3c6f */
            {8'h00}, /* 0x3c6e */
            {8'h00}, /* 0x3c6d */
            {8'h00}, /* 0x3c6c */
            {8'h00}, /* 0x3c6b */
            {8'h00}, /* 0x3c6a */
            {8'h00}, /* 0x3c69 */
            {8'h00}, /* 0x3c68 */
            {8'h00}, /* 0x3c67 */
            {8'h00}, /* 0x3c66 */
            {8'h00}, /* 0x3c65 */
            {8'h00}, /* 0x3c64 */
            {8'h00}, /* 0x3c63 */
            {8'h00}, /* 0x3c62 */
            {8'h00}, /* 0x3c61 */
            {8'h00}, /* 0x3c60 */
            {8'h00}, /* 0x3c5f */
            {8'h00}, /* 0x3c5e */
            {8'h00}, /* 0x3c5d */
            {8'h00}, /* 0x3c5c */
            {8'h00}, /* 0x3c5b */
            {8'h00}, /* 0x3c5a */
            {8'h00}, /* 0x3c59 */
            {8'h00}, /* 0x3c58 */
            {8'h00}, /* 0x3c57 */
            {8'h00}, /* 0x3c56 */
            {8'h00}, /* 0x3c55 */
            {8'h00}, /* 0x3c54 */
            {8'h00}, /* 0x3c53 */
            {8'h00}, /* 0x3c52 */
            {8'h00}, /* 0x3c51 */
            {8'h00}, /* 0x3c50 */
            {8'h00}, /* 0x3c4f */
            {8'h00}, /* 0x3c4e */
            {8'h00}, /* 0x3c4d */
            {8'h00}, /* 0x3c4c */
            {8'h00}, /* 0x3c4b */
            {8'h00}, /* 0x3c4a */
            {8'h00}, /* 0x3c49 */
            {8'h00}, /* 0x3c48 */
            {8'h00}, /* 0x3c47 */
            {8'h00}, /* 0x3c46 */
            {8'h00}, /* 0x3c45 */
            {8'h00}, /* 0x3c44 */
            {8'h00}, /* 0x3c43 */
            {8'h00}, /* 0x3c42 */
            {8'h00}, /* 0x3c41 */
            {8'h00}, /* 0x3c40 */
            {8'h00}, /* 0x3c3f */
            {8'h00}, /* 0x3c3e */
            {8'h00}, /* 0x3c3d */
            {8'h00}, /* 0x3c3c */
            {8'h00}, /* 0x3c3b */
            {8'h00}, /* 0x3c3a */
            {8'h00}, /* 0x3c39 */
            {8'h00}, /* 0x3c38 */
            {8'h00}, /* 0x3c37 */
            {8'h00}, /* 0x3c36 */
            {8'h00}, /* 0x3c35 */
            {8'h00}, /* 0x3c34 */
            {8'h00}, /* 0x3c33 */
            {8'h00}, /* 0x3c32 */
            {8'h00}, /* 0x3c31 */
            {8'h00}, /* 0x3c30 */
            {8'h00}, /* 0x3c2f */
            {8'h00}, /* 0x3c2e */
            {8'h00}, /* 0x3c2d */
            {8'h00}, /* 0x3c2c */
            {8'h00}, /* 0x3c2b */
            {8'h00}, /* 0x3c2a */
            {8'h00}, /* 0x3c29 */
            {8'h00}, /* 0x3c28 */
            {8'h00}, /* 0x3c27 */
            {8'h00}, /* 0x3c26 */
            {8'h00}, /* 0x3c25 */
            {8'h00}, /* 0x3c24 */
            {8'h00}, /* 0x3c23 */
            {8'h00}, /* 0x3c22 */
            {8'h00}, /* 0x3c21 */
            {8'h00}, /* 0x3c20 */
            {8'h00}, /* 0x3c1f */
            {8'h00}, /* 0x3c1e */
            {8'h00}, /* 0x3c1d */
            {8'h00}, /* 0x3c1c */
            {8'h00}, /* 0x3c1b */
            {8'h00}, /* 0x3c1a */
            {8'h00}, /* 0x3c19 */
            {8'h00}, /* 0x3c18 */
            {8'h00}, /* 0x3c17 */
            {8'h00}, /* 0x3c16 */
            {8'h00}, /* 0x3c15 */
            {8'h00}, /* 0x3c14 */
            {8'h00}, /* 0x3c13 */
            {8'h00}, /* 0x3c12 */
            {8'h00}, /* 0x3c11 */
            {8'h00}, /* 0x3c10 */
            {8'h00}, /* 0x3c0f */
            {8'h00}, /* 0x3c0e */
            {8'h00}, /* 0x3c0d */
            {8'h00}, /* 0x3c0c */
            {8'h00}, /* 0x3c0b */
            {8'h00}, /* 0x3c0a */
            {8'h00}, /* 0x3c09 */
            {8'h00}, /* 0x3c08 */
            {8'h00}, /* 0x3c07 */
            {8'h00}, /* 0x3c06 */
            {8'h00}, /* 0x3c05 */
            {8'h00}, /* 0x3c04 */
            {8'h00}, /* 0x3c03 */
            {8'h00}, /* 0x3c02 */
            {8'h00}, /* 0x3c01 */
            {8'h00}, /* 0x3c00 */
            {8'h00}, /* 0x3bff */
            {8'h00}, /* 0x3bfe */
            {8'h00}, /* 0x3bfd */
            {8'h00}, /* 0x3bfc */
            {8'h00}, /* 0x3bfb */
            {8'h00}, /* 0x3bfa */
            {8'h00}, /* 0x3bf9 */
            {8'h00}, /* 0x3bf8 */
            {8'h00}, /* 0x3bf7 */
            {8'h00}, /* 0x3bf6 */
            {8'h00}, /* 0x3bf5 */
            {8'h00}, /* 0x3bf4 */
            {8'h00}, /* 0x3bf3 */
            {8'h00}, /* 0x3bf2 */
            {8'h00}, /* 0x3bf1 */
            {8'h00}, /* 0x3bf0 */
            {8'h00}, /* 0x3bef */
            {8'h00}, /* 0x3bee */
            {8'h00}, /* 0x3bed */
            {8'h00}, /* 0x3bec */
            {8'h00}, /* 0x3beb */
            {8'h00}, /* 0x3bea */
            {8'h00}, /* 0x3be9 */
            {8'h00}, /* 0x3be8 */
            {8'h00}, /* 0x3be7 */
            {8'h00}, /* 0x3be6 */
            {8'h00}, /* 0x3be5 */
            {8'h00}, /* 0x3be4 */
            {8'h00}, /* 0x3be3 */
            {8'h00}, /* 0x3be2 */
            {8'h00}, /* 0x3be1 */
            {8'h00}, /* 0x3be0 */
            {8'h00}, /* 0x3bdf */
            {8'h00}, /* 0x3bde */
            {8'h00}, /* 0x3bdd */
            {8'h00}, /* 0x3bdc */
            {8'h00}, /* 0x3bdb */
            {8'h00}, /* 0x3bda */
            {8'h00}, /* 0x3bd9 */
            {8'h00}, /* 0x3bd8 */
            {8'h00}, /* 0x3bd7 */
            {8'h00}, /* 0x3bd6 */
            {8'h00}, /* 0x3bd5 */
            {8'h00}, /* 0x3bd4 */
            {8'h00}, /* 0x3bd3 */
            {8'h00}, /* 0x3bd2 */
            {8'h00}, /* 0x3bd1 */
            {8'h00}, /* 0x3bd0 */
            {8'h00}, /* 0x3bcf */
            {8'h00}, /* 0x3bce */
            {8'h00}, /* 0x3bcd */
            {8'h00}, /* 0x3bcc */
            {8'h00}, /* 0x3bcb */
            {8'h00}, /* 0x3bca */
            {8'h00}, /* 0x3bc9 */
            {8'h00}, /* 0x3bc8 */
            {8'h00}, /* 0x3bc7 */
            {8'h00}, /* 0x3bc6 */
            {8'h00}, /* 0x3bc5 */
            {8'h00}, /* 0x3bc4 */
            {8'h00}, /* 0x3bc3 */
            {8'h00}, /* 0x3bc2 */
            {8'h00}, /* 0x3bc1 */
            {8'h00}, /* 0x3bc0 */
            {8'h00}, /* 0x3bbf */
            {8'h00}, /* 0x3bbe */
            {8'h00}, /* 0x3bbd */
            {8'h00}, /* 0x3bbc */
            {8'h00}, /* 0x3bbb */
            {8'h00}, /* 0x3bba */
            {8'h00}, /* 0x3bb9 */
            {8'h00}, /* 0x3bb8 */
            {8'h00}, /* 0x3bb7 */
            {8'h00}, /* 0x3bb6 */
            {8'h00}, /* 0x3bb5 */
            {8'h00}, /* 0x3bb4 */
            {8'h00}, /* 0x3bb3 */
            {8'h00}, /* 0x3bb2 */
            {8'h00}, /* 0x3bb1 */
            {8'h00}, /* 0x3bb0 */
            {8'h00}, /* 0x3baf */
            {8'h00}, /* 0x3bae */
            {8'h00}, /* 0x3bad */
            {8'h00}, /* 0x3bac */
            {8'h00}, /* 0x3bab */
            {8'h00}, /* 0x3baa */
            {8'h00}, /* 0x3ba9 */
            {8'h00}, /* 0x3ba8 */
            {8'h00}, /* 0x3ba7 */
            {8'h00}, /* 0x3ba6 */
            {8'h00}, /* 0x3ba5 */
            {8'h00}, /* 0x3ba4 */
            {8'h00}, /* 0x3ba3 */
            {8'h00}, /* 0x3ba2 */
            {8'h00}, /* 0x3ba1 */
            {8'h00}, /* 0x3ba0 */
            {8'h00}, /* 0x3b9f */
            {8'h00}, /* 0x3b9e */
            {8'h00}, /* 0x3b9d */
            {8'h00}, /* 0x3b9c */
            {8'h00}, /* 0x3b9b */
            {8'h00}, /* 0x3b9a */
            {8'h00}, /* 0x3b99 */
            {8'h00}, /* 0x3b98 */
            {8'h00}, /* 0x3b97 */
            {8'h00}, /* 0x3b96 */
            {8'h00}, /* 0x3b95 */
            {8'h00}, /* 0x3b94 */
            {8'h00}, /* 0x3b93 */
            {8'h00}, /* 0x3b92 */
            {8'h00}, /* 0x3b91 */
            {8'h00}, /* 0x3b90 */
            {8'h00}, /* 0x3b8f */
            {8'h00}, /* 0x3b8e */
            {8'h00}, /* 0x3b8d */
            {8'h00}, /* 0x3b8c */
            {8'h00}, /* 0x3b8b */
            {8'h00}, /* 0x3b8a */
            {8'h00}, /* 0x3b89 */
            {8'h00}, /* 0x3b88 */
            {8'h00}, /* 0x3b87 */
            {8'h00}, /* 0x3b86 */
            {8'h00}, /* 0x3b85 */
            {8'h00}, /* 0x3b84 */
            {8'h00}, /* 0x3b83 */
            {8'h00}, /* 0x3b82 */
            {8'h00}, /* 0x3b81 */
            {8'h00}, /* 0x3b80 */
            {8'h00}, /* 0x3b7f */
            {8'h00}, /* 0x3b7e */
            {8'h00}, /* 0x3b7d */
            {8'h00}, /* 0x3b7c */
            {8'h00}, /* 0x3b7b */
            {8'h00}, /* 0x3b7a */
            {8'h00}, /* 0x3b79 */
            {8'h00}, /* 0x3b78 */
            {8'h00}, /* 0x3b77 */
            {8'h00}, /* 0x3b76 */
            {8'h00}, /* 0x3b75 */
            {8'h00}, /* 0x3b74 */
            {8'h00}, /* 0x3b73 */
            {8'h00}, /* 0x3b72 */
            {8'h00}, /* 0x3b71 */
            {8'h00}, /* 0x3b70 */
            {8'h00}, /* 0x3b6f */
            {8'h00}, /* 0x3b6e */
            {8'h00}, /* 0x3b6d */
            {8'h00}, /* 0x3b6c */
            {8'h00}, /* 0x3b6b */
            {8'h00}, /* 0x3b6a */
            {8'h00}, /* 0x3b69 */
            {8'h00}, /* 0x3b68 */
            {8'h00}, /* 0x3b67 */
            {8'h00}, /* 0x3b66 */
            {8'h00}, /* 0x3b65 */
            {8'h00}, /* 0x3b64 */
            {8'h00}, /* 0x3b63 */
            {8'h00}, /* 0x3b62 */
            {8'h00}, /* 0x3b61 */
            {8'h00}, /* 0x3b60 */
            {8'h00}, /* 0x3b5f */
            {8'h00}, /* 0x3b5e */
            {8'h00}, /* 0x3b5d */
            {8'h00}, /* 0x3b5c */
            {8'h00}, /* 0x3b5b */
            {8'h00}, /* 0x3b5a */
            {8'h00}, /* 0x3b59 */
            {8'h00}, /* 0x3b58 */
            {8'h00}, /* 0x3b57 */
            {8'h00}, /* 0x3b56 */
            {8'h00}, /* 0x3b55 */
            {8'h00}, /* 0x3b54 */
            {8'h00}, /* 0x3b53 */
            {8'h00}, /* 0x3b52 */
            {8'h00}, /* 0x3b51 */
            {8'h00}, /* 0x3b50 */
            {8'h00}, /* 0x3b4f */
            {8'h00}, /* 0x3b4e */
            {8'h00}, /* 0x3b4d */
            {8'h00}, /* 0x3b4c */
            {8'h00}, /* 0x3b4b */
            {8'h00}, /* 0x3b4a */
            {8'h00}, /* 0x3b49 */
            {8'h00}, /* 0x3b48 */
            {8'h00}, /* 0x3b47 */
            {8'h00}, /* 0x3b46 */
            {8'h00}, /* 0x3b45 */
            {8'h00}, /* 0x3b44 */
            {8'h00}, /* 0x3b43 */
            {8'h00}, /* 0x3b42 */
            {8'h00}, /* 0x3b41 */
            {8'h00}, /* 0x3b40 */
            {8'h00}, /* 0x3b3f */
            {8'h00}, /* 0x3b3e */
            {8'h00}, /* 0x3b3d */
            {8'h00}, /* 0x3b3c */
            {8'h00}, /* 0x3b3b */
            {8'h00}, /* 0x3b3a */
            {8'h00}, /* 0x3b39 */
            {8'h00}, /* 0x3b38 */
            {8'h00}, /* 0x3b37 */
            {8'h00}, /* 0x3b36 */
            {8'h00}, /* 0x3b35 */
            {8'h00}, /* 0x3b34 */
            {8'h00}, /* 0x3b33 */
            {8'h00}, /* 0x3b32 */
            {8'h00}, /* 0x3b31 */
            {8'h00}, /* 0x3b30 */
            {8'h00}, /* 0x3b2f */
            {8'h00}, /* 0x3b2e */
            {8'h00}, /* 0x3b2d */
            {8'h00}, /* 0x3b2c */
            {8'h00}, /* 0x3b2b */
            {8'h00}, /* 0x3b2a */
            {8'h00}, /* 0x3b29 */
            {8'h00}, /* 0x3b28 */
            {8'h00}, /* 0x3b27 */
            {8'h00}, /* 0x3b26 */
            {8'h00}, /* 0x3b25 */
            {8'h00}, /* 0x3b24 */
            {8'h00}, /* 0x3b23 */
            {8'h00}, /* 0x3b22 */
            {8'h00}, /* 0x3b21 */
            {8'h00}, /* 0x3b20 */
            {8'h00}, /* 0x3b1f */
            {8'h00}, /* 0x3b1e */
            {8'h00}, /* 0x3b1d */
            {8'h00}, /* 0x3b1c */
            {8'h00}, /* 0x3b1b */
            {8'h00}, /* 0x3b1a */
            {8'h00}, /* 0x3b19 */
            {8'h00}, /* 0x3b18 */
            {8'h00}, /* 0x3b17 */
            {8'h00}, /* 0x3b16 */
            {8'h00}, /* 0x3b15 */
            {8'h00}, /* 0x3b14 */
            {8'h00}, /* 0x3b13 */
            {8'h00}, /* 0x3b12 */
            {8'h00}, /* 0x3b11 */
            {8'h00}, /* 0x3b10 */
            {8'h00}, /* 0x3b0f */
            {8'h00}, /* 0x3b0e */
            {8'h00}, /* 0x3b0d */
            {8'h00}, /* 0x3b0c */
            {8'h00}, /* 0x3b0b */
            {8'h00}, /* 0x3b0a */
            {8'h00}, /* 0x3b09 */
            {8'h00}, /* 0x3b08 */
            {8'h00}, /* 0x3b07 */
            {8'h00}, /* 0x3b06 */
            {8'h00}, /* 0x3b05 */
            {8'h00}, /* 0x3b04 */
            {8'h00}, /* 0x3b03 */
            {8'h00}, /* 0x3b02 */
            {8'h00}, /* 0x3b01 */
            {8'h00}, /* 0x3b00 */
            {8'h00}, /* 0x3aff */
            {8'h00}, /* 0x3afe */
            {8'h00}, /* 0x3afd */
            {8'h00}, /* 0x3afc */
            {8'h00}, /* 0x3afb */
            {8'h00}, /* 0x3afa */
            {8'h00}, /* 0x3af9 */
            {8'h00}, /* 0x3af8 */
            {8'h00}, /* 0x3af7 */
            {8'h00}, /* 0x3af6 */
            {8'h00}, /* 0x3af5 */
            {8'h00}, /* 0x3af4 */
            {8'h00}, /* 0x3af3 */
            {8'h00}, /* 0x3af2 */
            {8'h00}, /* 0x3af1 */
            {8'h00}, /* 0x3af0 */
            {8'h00}, /* 0x3aef */
            {8'h00}, /* 0x3aee */
            {8'h00}, /* 0x3aed */
            {8'h00}, /* 0x3aec */
            {8'h00}, /* 0x3aeb */
            {8'h00}, /* 0x3aea */
            {8'h00}, /* 0x3ae9 */
            {8'h00}, /* 0x3ae8 */
            {8'h00}, /* 0x3ae7 */
            {8'h00}, /* 0x3ae6 */
            {8'h00}, /* 0x3ae5 */
            {8'h00}, /* 0x3ae4 */
            {8'h00}, /* 0x3ae3 */
            {8'h00}, /* 0x3ae2 */
            {8'h00}, /* 0x3ae1 */
            {8'h00}, /* 0x3ae0 */
            {8'h00}, /* 0x3adf */
            {8'h00}, /* 0x3ade */
            {8'h00}, /* 0x3add */
            {8'h00}, /* 0x3adc */
            {8'h00}, /* 0x3adb */
            {8'h00}, /* 0x3ada */
            {8'h00}, /* 0x3ad9 */
            {8'h00}, /* 0x3ad8 */
            {8'h00}, /* 0x3ad7 */
            {8'h00}, /* 0x3ad6 */
            {8'h00}, /* 0x3ad5 */
            {8'h00}, /* 0x3ad4 */
            {8'h00}, /* 0x3ad3 */
            {8'h00}, /* 0x3ad2 */
            {8'h00}, /* 0x3ad1 */
            {8'h00}, /* 0x3ad0 */
            {8'h00}, /* 0x3acf */
            {8'h00}, /* 0x3ace */
            {8'h00}, /* 0x3acd */
            {8'h00}, /* 0x3acc */
            {8'h00}, /* 0x3acb */
            {8'h00}, /* 0x3aca */
            {8'h00}, /* 0x3ac9 */
            {8'h00}, /* 0x3ac8 */
            {8'h00}, /* 0x3ac7 */
            {8'h00}, /* 0x3ac6 */
            {8'h00}, /* 0x3ac5 */
            {8'h00}, /* 0x3ac4 */
            {8'h00}, /* 0x3ac3 */
            {8'h00}, /* 0x3ac2 */
            {8'h00}, /* 0x3ac1 */
            {8'h00}, /* 0x3ac0 */
            {8'h00}, /* 0x3abf */
            {8'h00}, /* 0x3abe */
            {8'h00}, /* 0x3abd */
            {8'h00}, /* 0x3abc */
            {8'h00}, /* 0x3abb */
            {8'h00}, /* 0x3aba */
            {8'h00}, /* 0x3ab9 */
            {8'h00}, /* 0x3ab8 */
            {8'h00}, /* 0x3ab7 */
            {8'h00}, /* 0x3ab6 */
            {8'h00}, /* 0x3ab5 */
            {8'h00}, /* 0x3ab4 */
            {8'h00}, /* 0x3ab3 */
            {8'h00}, /* 0x3ab2 */
            {8'h00}, /* 0x3ab1 */
            {8'h00}, /* 0x3ab0 */
            {8'h00}, /* 0x3aaf */
            {8'h00}, /* 0x3aae */
            {8'h00}, /* 0x3aad */
            {8'h00}, /* 0x3aac */
            {8'h00}, /* 0x3aab */
            {8'h00}, /* 0x3aaa */
            {8'h00}, /* 0x3aa9 */
            {8'h00}, /* 0x3aa8 */
            {8'h00}, /* 0x3aa7 */
            {8'h00}, /* 0x3aa6 */
            {8'h00}, /* 0x3aa5 */
            {8'h00}, /* 0x3aa4 */
            {8'h00}, /* 0x3aa3 */
            {8'h00}, /* 0x3aa2 */
            {8'h00}, /* 0x3aa1 */
            {8'h00}, /* 0x3aa0 */
            {8'h00}, /* 0x3a9f */
            {8'h00}, /* 0x3a9e */
            {8'h00}, /* 0x3a9d */
            {8'h00}, /* 0x3a9c */
            {8'h00}, /* 0x3a9b */
            {8'h00}, /* 0x3a9a */
            {8'h00}, /* 0x3a99 */
            {8'h00}, /* 0x3a98 */
            {8'h00}, /* 0x3a97 */
            {8'h00}, /* 0x3a96 */
            {8'h00}, /* 0x3a95 */
            {8'h00}, /* 0x3a94 */
            {8'h00}, /* 0x3a93 */
            {8'h00}, /* 0x3a92 */
            {8'h00}, /* 0x3a91 */
            {8'h00}, /* 0x3a90 */
            {8'h00}, /* 0x3a8f */
            {8'h00}, /* 0x3a8e */
            {8'h00}, /* 0x3a8d */
            {8'h00}, /* 0x3a8c */
            {8'h00}, /* 0x3a8b */
            {8'h00}, /* 0x3a8a */
            {8'h00}, /* 0x3a89 */
            {8'h00}, /* 0x3a88 */
            {8'h00}, /* 0x3a87 */
            {8'h00}, /* 0x3a86 */
            {8'h00}, /* 0x3a85 */
            {8'h00}, /* 0x3a84 */
            {8'h00}, /* 0x3a83 */
            {8'h00}, /* 0x3a82 */
            {8'h00}, /* 0x3a81 */
            {8'h00}, /* 0x3a80 */
            {8'h00}, /* 0x3a7f */
            {8'h00}, /* 0x3a7e */
            {8'h00}, /* 0x3a7d */
            {8'h00}, /* 0x3a7c */
            {8'h00}, /* 0x3a7b */
            {8'h00}, /* 0x3a7a */
            {8'h00}, /* 0x3a79 */
            {8'h00}, /* 0x3a78 */
            {8'h00}, /* 0x3a77 */
            {8'h00}, /* 0x3a76 */
            {8'h00}, /* 0x3a75 */
            {8'h00}, /* 0x3a74 */
            {8'h00}, /* 0x3a73 */
            {8'h00}, /* 0x3a72 */
            {8'h00}, /* 0x3a71 */
            {8'h00}, /* 0x3a70 */
            {8'h00}, /* 0x3a6f */
            {8'h00}, /* 0x3a6e */
            {8'h00}, /* 0x3a6d */
            {8'h00}, /* 0x3a6c */
            {8'h00}, /* 0x3a6b */
            {8'h00}, /* 0x3a6a */
            {8'h00}, /* 0x3a69 */
            {8'h00}, /* 0x3a68 */
            {8'h00}, /* 0x3a67 */
            {8'h00}, /* 0x3a66 */
            {8'h00}, /* 0x3a65 */
            {8'h00}, /* 0x3a64 */
            {8'h00}, /* 0x3a63 */
            {8'h00}, /* 0x3a62 */
            {8'h00}, /* 0x3a61 */
            {8'h00}, /* 0x3a60 */
            {8'h00}, /* 0x3a5f */
            {8'h00}, /* 0x3a5e */
            {8'h00}, /* 0x3a5d */
            {8'h00}, /* 0x3a5c */
            {8'h00}, /* 0x3a5b */
            {8'h00}, /* 0x3a5a */
            {8'h00}, /* 0x3a59 */
            {8'h00}, /* 0x3a58 */
            {8'h00}, /* 0x3a57 */
            {8'h00}, /* 0x3a56 */
            {8'h00}, /* 0x3a55 */
            {8'h00}, /* 0x3a54 */
            {8'h00}, /* 0x3a53 */
            {8'h00}, /* 0x3a52 */
            {8'h00}, /* 0x3a51 */
            {8'h00}, /* 0x3a50 */
            {8'h00}, /* 0x3a4f */
            {8'h00}, /* 0x3a4e */
            {8'h00}, /* 0x3a4d */
            {8'h00}, /* 0x3a4c */
            {8'h00}, /* 0x3a4b */
            {8'h00}, /* 0x3a4a */
            {8'h00}, /* 0x3a49 */
            {8'h00}, /* 0x3a48 */
            {8'h00}, /* 0x3a47 */
            {8'h00}, /* 0x3a46 */
            {8'h00}, /* 0x3a45 */
            {8'h00}, /* 0x3a44 */
            {8'h00}, /* 0x3a43 */
            {8'h00}, /* 0x3a42 */
            {8'h00}, /* 0x3a41 */
            {8'h00}, /* 0x3a40 */
            {8'h00}, /* 0x3a3f */
            {8'h00}, /* 0x3a3e */
            {8'h00}, /* 0x3a3d */
            {8'h00}, /* 0x3a3c */
            {8'h00}, /* 0x3a3b */
            {8'h00}, /* 0x3a3a */
            {8'h00}, /* 0x3a39 */
            {8'h00}, /* 0x3a38 */
            {8'h00}, /* 0x3a37 */
            {8'h00}, /* 0x3a36 */
            {8'h00}, /* 0x3a35 */
            {8'h00}, /* 0x3a34 */
            {8'h00}, /* 0x3a33 */
            {8'h00}, /* 0x3a32 */
            {8'h00}, /* 0x3a31 */
            {8'h00}, /* 0x3a30 */
            {8'h00}, /* 0x3a2f */
            {8'h00}, /* 0x3a2e */
            {8'h00}, /* 0x3a2d */
            {8'h00}, /* 0x3a2c */
            {8'h00}, /* 0x3a2b */
            {8'h00}, /* 0x3a2a */
            {8'h00}, /* 0x3a29 */
            {8'h00}, /* 0x3a28 */
            {8'h00}, /* 0x3a27 */
            {8'h00}, /* 0x3a26 */
            {8'h00}, /* 0x3a25 */
            {8'h00}, /* 0x3a24 */
            {8'h00}, /* 0x3a23 */
            {8'h00}, /* 0x3a22 */
            {8'h00}, /* 0x3a21 */
            {8'h00}, /* 0x3a20 */
            {8'h00}, /* 0x3a1f */
            {8'h00}, /* 0x3a1e */
            {8'h00}, /* 0x3a1d */
            {8'h00}, /* 0x3a1c */
            {8'h00}, /* 0x3a1b */
            {8'h00}, /* 0x3a1a */
            {8'h00}, /* 0x3a19 */
            {8'h00}, /* 0x3a18 */
            {8'h00}, /* 0x3a17 */
            {8'h00}, /* 0x3a16 */
            {8'h00}, /* 0x3a15 */
            {8'h00}, /* 0x3a14 */
            {8'h00}, /* 0x3a13 */
            {8'h00}, /* 0x3a12 */
            {8'h00}, /* 0x3a11 */
            {8'h00}, /* 0x3a10 */
            {8'h00}, /* 0x3a0f */
            {8'h00}, /* 0x3a0e */
            {8'h00}, /* 0x3a0d */
            {8'h00}, /* 0x3a0c */
            {8'h00}, /* 0x3a0b */
            {8'h00}, /* 0x3a0a */
            {8'h00}, /* 0x3a09 */
            {8'h00}, /* 0x3a08 */
            {8'h00}, /* 0x3a07 */
            {8'h00}, /* 0x3a06 */
            {8'h00}, /* 0x3a05 */
            {8'h00}, /* 0x3a04 */
            {8'h00}, /* 0x3a03 */
            {8'h00}, /* 0x3a02 */
            {8'h00}, /* 0x3a01 */
            {8'h00}, /* 0x3a00 */
            {8'h00}, /* 0x39ff */
            {8'h00}, /* 0x39fe */
            {8'h00}, /* 0x39fd */
            {8'h00}, /* 0x39fc */
            {8'h00}, /* 0x39fb */
            {8'h00}, /* 0x39fa */
            {8'h00}, /* 0x39f9 */
            {8'h00}, /* 0x39f8 */
            {8'h00}, /* 0x39f7 */
            {8'h00}, /* 0x39f6 */
            {8'h00}, /* 0x39f5 */
            {8'h00}, /* 0x39f4 */
            {8'h00}, /* 0x39f3 */
            {8'h00}, /* 0x39f2 */
            {8'h00}, /* 0x39f1 */
            {8'h00}, /* 0x39f0 */
            {8'h00}, /* 0x39ef */
            {8'h00}, /* 0x39ee */
            {8'h00}, /* 0x39ed */
            {8'h00}, /* 0x39ec */
            {8'h00}, /* 0x39eb */
            {8'h00}, /* 0x39ea */
            {8'h00}, /* 0x39e9 */
            {8'h00}, /* 0x39e8 */
            {8'h00}, /* 0x39e7 */
            {8'h00}, /* 0x39e6 */
            {8'h00}, /* 0x39e5 */
            {8'h00}, /* 0x39e4 */
            {8'h00}, /* 0x39e3 */
            {8'h00}, /* 0x39e2 */
            {8'h00}, /* 0x39e1 */
            {8'h00}, /* 0x39e0 */
            {8'h00}, /* 0x39df */
            {8'h00}, /* 0x39de */
            {8'h00}, /* 0x39dd */
            {8'h00}, /* 0x39dc */
            {8'h00}, /* 0x39db */
            {8'h00}, /* 0x39da */
            {8'h00}, /* 0x39d9 */
            {8'h00}, /* 0x39d8 */
            {8'h00}, /* 0x39d7 */
            {8'h00}, /* 0x39d6 */
            {8'h00}, /* 0x39d5 */
            {8'h00}, /* 0x39d4 */
            {8'h00}, /* 0x39d3 */
            {8'h00}, /* 0x39d2 */
            {8'h00}, /* 0x39d1 */
            {8'h00}, /* 0x39d0 */
            {8'h00}, /* 0x39cf */
            {8'h00}, /* 0x39ce */
            {8'h00}, /* 0x39cd */
            {8'h00}, /* 0x39cc */
            {8'h00}, /* 0x39cb */
            {8'h00}, /* 0x39ca */
            {8'h00}, /* 0x39c9 */
            {8'h00}, /* 0x39c8 */
            {8'h00}, /* 0x39c7 */
            {8'h00}, /* 0x39c6 */
            {8'h00}, /* 0x39c5 */
            {8'h00}, /* 0x39c4 */
            {8'h00}, /* 0x39c3 */
            {8'h00}, /* 0x39c2 */
            {8'h00}, /* 0x39c1 */
            {8'h00}, /* 0x39c0 */
            {8'h00}, /* 0x39bf */
            {8'h00}, /* 0x39be */
            {8'h00}, /* 0x39bd */
            {8'h00}, /* 0x39bc */
            {8'h00}, /* 0x39bb */
            {8'h00}, /* 0x39ba */
            {8'h00}, /* 0x39b9 */
            {8'h00}, /* 0x39b8 */
            {8'h00}, /* 0x39b7 */
            {8'h00}, /* 0x39b6 */
            {8'h00}, /* 0x39b5 */
            {8'h00}, /* 0x39b4 */
            {8'h00}, /* 0x39b3 */
            {8'h00}, /* 0x39b2 */
            {8'h00}, /* 0x39b1 */
            {8'h00}, /* 0x39b0 */
            {8'h00}, /* 0x39af */
            {8'h00}, /* 0x39ae */
            {8'h00}, /* 0x39ad */
            {8'h00}, /* 0x39ac */
            {8'h00}, /* 0x39ab */
            {8'h00}, /* 0x39aa */
            {8'h00}, /* 0x39a9 */
            {8'h00}, /* 0x39a8 */
            {8'h00}, /* 0x39a7 */
            {8'h00}, /* 0x39a6 */
            {8'h00}, /* 0x39a5 */
            {8'h00}, /* 0x39a4 */
            {8'h00}, /* 0x39a3 */
            {8'h00}, /* 0x39a2 */
            {8'h00}, /* 0x39a1 */
            {8'h00}, /* 0x39a0 */
            {8'h00}, /* 0x399f */
            {8'h00}, /* 0x399e */
            {8'h00}, /* 0x399d */
            {8'h00}, /* 0x399c */
            {8'h00}, /* 0x399b */
            {8'h00}, /* 0x399a */
            {8'h00}, /* 0x3999 */
            {8'h00}, /* 0x3998 */
            {8'h00}, /* 0x3997 */
            {8'h00}, /* 0x3996 */
            {8'h00}, /* 0x3995 */
            {8'h00}, /* 0x3994 */
            {8'h00}, /* 0x3993 */
            {8'h00}, /* 0x3992 */
            {8'h00}, /* 0x3991 */
            {8'h00}, /* 0x3990 */
            {8'h00}, /* 0x398f */
            {8'h00}, /* 0x398e */
            {8'h00}, /* 0x398d */
            {8'h00}, /* 0x398c */
            {8'h00}, /* 0x398b */
            {8'h00}, /* 0x398a */
            {8'h00}, /* 0x3989 */
            {8'h00}, /* 0x3988 */
            {8'h00}, /* 0x3987 */
            {8'h00}, /* 0x3986 */
            {8'h00}, /* 0x3985 */
            {8'h00}, /* 0x3984 */
            {8'h00}, /* 0x3983 */
            {8'h00}, /* 0x3982 */
            {8'h00}, /* 0x3981 */
            {8'h00}, /* 0x3980 */
            {8'h00}, /* 0x397f */
            {8'h00}, /* 0x397e */
            {8'h00}, /* 0x397d */
            {8'h00}, /* 0x397c */
            {8'h00}, /* 0x397b */
            {8'h00}, /* 0x397a */
            {8'h00}, /* 0x3979 */
            {8'h00}, /* 0x3978 */
            {8'h00}, /* 0x3977 */
            {8'h00}, /* 0x3976 */
            {8'h00}, /* 0x3975 */
            {8'h00}, /* 0x3974 */
            {8'h00}, /* 0x3973 */
            {8'h00}, /* 0x3972 */
            {8'h00}, /* 0x3971 */
            {8'h00}, /* 0x3970 */
            {8'h00}, /* 0x396f */
            {8'h00}, /* 0x396e */
            {8'h00}, /* 0x396d */
            {8'h00}, /* 0x396c */
            {8'h00}, /* 0x396b */
            {8'h00}, /* 0x396a */
            {8'h00}, /* 0x3969 */
            {8'h00}, /* 0x3968 */
            {8'h00}, /* 0x3967 */
            {8'h00}, /* 0x3966 */
            {8'h00}, /* 0x3965 */
            {8'h00}, /* 0x3964 */
            {8'h00}, /* 0x3963 */
            {8'h00}, /* 0x3962 */
            {8'h00}, /* 0x3961 */
            {8'h00}, /* 0x3960 */
            {8'h00}, /* 0x395f */
            {8'h00}, /* 0x395e */
            {8'h00}, /* 0x395d */
            {8'h00}, /* 0x395c */
            {8'h00}, /* 0x395b */
            {8'h00}, /* 0x395a */
            {8'h00}, /* 0x3959 */
            {8'h00}, /* 0x3958 */
            {8'h00}, /* 0x3957 */
            {8'h00}, /* 0x3956 */
            {8'h00}, /* 0x3955 */
            {8'h00}, /* 0x3954 */
            {8'h00}, /* 0x3953 */
            {8'h00}, /* 0x3952 */
            {8'h00}, /* 0x3951 */
            {8'h00}, /* 0x3950 */
            {8'h00}, /* 0x394f */
            {8'h00}, /* 0x394e */
            {8'h00}, /* 0x394d */
            {8'h00}, /* 0x394c */
            {8'h00}, /* 0x394b */
            {8'h00}, /* 0x394a */
            {8'h00}, /* 0x3949 */
            {8'h00}, /* 0x3948 */
            {8'h00}, /* 0x3947 */
            {8'h00}, /* 0x3946 */
            {8'h00}, /* 0x3945 */
            {8'h00}, /* 0x3944 */
            {8'h00}, /* 0x3943 */
            {8'h00}, /* 0x3942 */
            {8'h00}, /* 0x3941 */
            {8'h00}, /* 0x3940 */
            {8'h00}, /* 0x393f */
            {8'h00}, /* 0x393e */
            {8'h00}, /* 0x393d */
            {8'h00}, /* 0x393c */
            {8'h00}, /* 0x393b */
            {8'h00}, /* 0x393a */
            {8'h00}, /* 0x3939 */
            {8'h00}, /* 0x3938 */
            {8'h00}, /* 0x3937 */
            {8'h00}, /* 0x3936 */
            {8'h00}, /* 0x3935 */
            {8'h00}, /* 0x3934 */
            {8'h00}, /* 0x3933 */
            {8'h00}, /* 0x3932 */
            {8'h00}, /* 0x3931 */
            {8'h00}, /* 0x3930 */
            {8'h00}, /* 0x392f */
            {8'h00}, /* 0x392e */
            {8'h00}, /* 0x392d */
            {8'h00}, /* 0x392c */
            {8'h00}, /* 0x392b */
            {8'h00}, /* 0x392a */
            {8'h00}, /* 0x3929 */
            {8'h00}, /* 0x3928 */
            {8'h00}, /* 0x3927 */
            {8'h00}, /* 0x3926 */
            {8'h00}, /* 0x3925 */
            {8'h00}, /* 0x3924 */
            {8'h00}, /* 0x3923 */
            {8'h00}, /* 0x3922 */
            {8'h00}, /* 0x3921 */
            {8'h00}, /* 0x3920 */
            {8'h00}, /* 0x391f */
            {8'h00}, /* 0x391e */
            {8'h00}, /* 0x391d */
            {8'h00}, /* 0x391c */
            {8'h00}, /* 0x391b */
            {8'h00}, /* 0x391a */
            {8'h00}, /* 0x3919 */
            {8'h00}, /* 0x3918 */
            {8'h00}, /* 0x3917 */
            {8'h00}, /* 0x3916 */
            {8'h00}, /* 0x3915 */
            {8'h00}, /* 0x3914 */
            {8'h00}, /* 0x3913 */
            {8'h00}, /* 0x3912 */
            {8'h00}, /* 0x3911 */
            {8'h00}, /* 0x3910 */
            {8'h00}, /* 0x390f */
            {8'h00}, /* 0x390e */
            {8'h00}, /* 0x390d */
            {8'h00}, /* 0x390c */
            {8'h00}, /* 0x390b */
            {8'h00}, /* 0x390a */
            {8'h00}, /* 0x3909 */
            {8'h00}, /* 0x3908 */
            {8'h00}, /* 0x3907 */
            {8'h00}, /* 0x3906 */
            {8'h00}, /* 0x3905 */
            {8'h00}, /* 0x3904 */
            {8'h00}, /* 0x3903 */
            {8'h00}, /* 0x3902 */
            {8'h00}, /* 0x3901 */
            {8'h00}, /* 0x3900 */
            {8'h00}, /* 0x38ff */
            {8'h00}, /* 0x38fe */
            {8'h00}, /* 0x38fd */
            {8'h00}, /* 0x38fc */
            {8'h00}, /* 0x38fb */
            {8'h00}, /* 0x38fa */
            {8'h00}, /* 0x38f9 */
            {8'h00}, /* 0x38f8 */
            {8'h00}, /* 0x38f7 */
            {8'h00}, /* 0x38f6 */
            {8'h00}, /* 0x38f5 */
            {8'h00}, /* 0x38f4 */
            {8'h00}, /* 0x38f3 */
            {8'h00}, /* 0x38f2 */
            {8'h00}, /* 0x38f1 */
            {8'h00}, /* 0x38f0 */
            {8'h00}, /* 0x38ef */
            {8'h00}, /* 0x38ee */
            {8'h00}, /* 0x38ed */
            {8'h00}, /* 0x38ec */
            {8'h00}, /* 0x38eb */
            {8'h00}, /* 0x38ea */
            {8'h00}, /* 0x38e9 */
            {8'h00}, /* 0x38e8 */
            {8'h00}, /* 0x38e7 */
            {8'h00}, /* 0x38e6 */
            {8'h00}, /* 0x38e5 */
            {8'h00}, /* 0x38e4 */
            {8'h00}, /* 0x38e3 */
            {8'h00}, /* 0x38e2 */
            {8'h00}, /* 0x38e1 */
            {8'h00}, /* 0x38e0 */
            {8'h00}, /* 0x38df */
            {8'h00}, /* 0x38de */
            {8'h00}, /* 0x38dd */
            {8'h00}, /* 0x38dc */
            {8'h00}, /* 0x38db */
            {8'h00}, /* 0x38da */
            {8'h00}, /* 0x38d9 */
            {8'h00}, /* 0x38d8 */
            {8'h00}, /* 0x38d7 */
            {8'h00}, /* 0x38d6 */
            {8'h00}, /* 0x38d5 */
            {8'h00}, /* 0x38d4 */
            {8'h00}, /* 0x38d3 */
            {8'h00}, /* 0x38d2 */
            {8'h00}, /* 0x38d1 */
            {8'h00}, /* 0x38d0 */
            {8'h00}, /* 0x38cf */
            {8'h00}, /* 0x38ce */
            {8'h00}, /* 0x38cd */
            {8'h00}, /* 0x38cc */
            {8'h00}, /* 0x38cb */
            {8'h00}, /* 0x38ca */
            {8'h00}, /* 0x38c9 */
            {8'h00}, /* 0x38c8 */
            {8'h00}, /* 0x38c7 */
            {8'h00}, /* 0x38c6 */
            {8'h00}, /* 0x38c5 */
            {8'h00}, /* 0x38c4 */
            {8'h00}, /* 0x38c3 */
            {8'h00}, /* 0x38c2 */
            {8'h00}, /* 0x38c1 */
            {8'h00}, /* 0x38c0 */
            {8'h00}, /* 0x38bf */
            {8'h00}, /* 0x38be */
            {8'h00}, /* 0x38bd */
            {8'h00}, /* 0x38bc */
            {8'h00}, /* 0x38bb */
            {8'h00}, /* 0x38ba */
            {8'h00}, /* 0x38b9 */
            {8'h00}, /* 0x38b8 */
            {8'h00}, /* 0x38b7 */
            {8'h00}, /* 0x38b6 */
            {8'h00}, /* 0x38b5 */
            {8'h00}, /* 0x38b4 */
            {8'h00}, /* 0x38b3 */
            {8'h00}, /* 0x38b2 */
            {8'h00}, /* 0x38b1 */
            {8'h00}, /* 0x38b0 */
            {8'h00}, /* 0x38af */
            {8'h00}, /* 0x38ae */
            {8'h00}, /* 0x38ad */
            {8'h00}, /* 0x38ac */
            {8'h00}, /* 0x38ab */
            {8'h00}, /* 0x38aa */
            {8'h00}, /* 0x38a9 */
            {8'h00}, /* 0x38a8 */
            {8'h00}, /* 0x38a7 */
            {8'h00}, /* 0x38a6 */
            {8'h00}, /* 0x38a5 */
            {8'h00}, /* 0x38a4 */
            {8'h00}, /* 0x38a3 */
            {8'h00}, /* 0x38a2 */
            {8'h00}, /* 0x38a1 */
            {8'h00}, /* 0x38a0 */
            {8'h00}, /* 0x389f */
            {8'h00}, /* 0x389e */
            {8'h00}, /* 0x389d */
            {8'h00}, /* 0x389c */
            {8'h00}, /* 0x389b */
            {8'h00}, /* 0x389a */
            {8'h00}, /* 0x3899 */
            {8'h00}, /* 0x3898 */
            {8'h00}, /* 0x3897 */
            {8'h00}, /* 0x3896 */
            {8'h00}, /* 0x3895 */
            {8'h00}, /* 0x3894 */
            {8'h00}, /* 0x3893 */
            {8'h00}, /* 0x3892 */
            {8'h00}, /* 0x3891 */
            {8'h00}, /* 0x3890 */
            {8'h00}, /* 0x388f */
            {8'h00}, /* 0x388e */
            {8'h00}, /* 0x388d */
            {8'h00}, /* 0x388c */
            {8'h00}, /* 0x388b */
            {8'h00}, /* 0x388a */
            {8'h00}, /* 0x3889 */
            {8'h00}, /* 0x3888 */
            {8'h00}, /* 0x3887 */
            {8'h00}, /* 0x3886 */
            {8'h00}, /* 0x3885 */
            {8'h00}, /* 0x3884 */
            {8'h00}, /* 0x3883 */
            {8'h00}, /* 0x3882 */
            {8'h00}, /* 0x3881 */
            {8'h00}, /* 0x3880 */
            {8'h00}, /* 0x387f */
            {8'h00}, /* 0x387e */
            {8'h00}, /* 0x387d */
            {8'h00}, /* 0x387c */
            {8'h00}, /* 0x387b */
            {8'h00}, /* 0x387a */
            {8'h00}, /* 0x3879 */
            {8'h00}, /* 0x3878 */
            {8'h00}, /* 0x3877 */
            {8'h00}, /* 0x3876 */
            {8'h00}, /* 0x3875 */
            {8'h00}, /* 0x3874 */
            {8'h00}, /* 0x3873 */
            {8'h00}, /* 0x3872 */
            {8'h00}, /* 0x3871 */
            {8'h00}, /* 0x3870 */
            {8'h00}, /* 0x386f */
            {8'h00}, /* 0x386e */
            {8'h00}, /* 0x386d */
            {8'h00}, /* 0x386c */
            {8'h00}, /* 0x386b */
            {8'h00}, /* 0x386a */
            {8'h00}, /* 0x3869 */
            {8'h00}, /* 0x3868 */
            {8'h00}, /* 0x3867 */
            {8'h00}, /* 0x3866 */
            {8'h00}, /* 0x3865 */
            {8'h00}, /* 0x3864 */
            {8'h00}, /* 0x3863 */
            {8'h00}, /* 0x3862 */
            {8'h00}, /* 0x3861 */
            {8'h00}, /* 0x3860 */
            {8'h00}, /* 0x385f */
            {8'h00}, /* 0x385e */
            {8'h00}, /* 0x385d */
            {8'h00}, /* 0x385c */
            {8'h00}, /* 0x385b */
            {8'h00}, /* 0x385a */
            {8'h00}, /* 0x3859 */
            {8'h00}, /* 0x3858 */
            {8'h00}, /* 0x3857 */
            {8'h00}, /* 0x3856 */
            {8'h00}, /* 0x3855 */
            {8'h00}, /* 0x3854 */
            {8'h00}, /* 0x3853 */
            {8'h00}, /* 0x3852 */
            {8'h00}, /* 0x3851 */
            {8'h00}, /* 0x3850 */
            {8'h00}, /* 0x384f */
            {8'h00}, /* 0x384e */
            {8'h00}, /* 0x384d */
            {8'h00}, /* 0x384c */
            {8'h00}, /* 0x384b */
            {8'h00}, /* 0x384a */
            {8'h00}, /* 0x3849 */
            {8'h00}, /* 0x3848 */
            {8'h00}, /* 0x3847 */
            {8'h00}, /* 0x3846 */
            {8'h00}, /* 0x3845 */
            {8'h00}, /* 0x3844 */
            {8'h00}, /* 0x3843 */
            {8'h00}, /* 0x3842 */
            {8'h00}, /* 0x3841 */
            {8'h00}, /* 0x3840 */
            {8'h00}, /* 0x383f */
            {8'h00}, /* 0x383e */
            {8'h00}, /* 0x383d */
            {8'h00}, /* 0x383c */
            {8'h00}, /* 0x383b */
            {8'h00}, /* 0x383a */
            {8'h00}, /* 0x3839 */
            {8'h00}, /* 0x3838 */
            {8'h00}, /* 0x3837 */
            {8'h00}, /* 0x3836 */
            {8'h00}, /* 0x3835 */
            {8'h00}, /* 0x3834 */
            {8'h00}, /* 0x3833 */
            {8'h00}, /* 0x3832 */
            {8'h00}, /* 0x3831 */
            {8'h00}, /* 0x3830 */
            {8'h00}, /* 0x382f */
            {8'h00}, /* 0x382e */
            {8'h00}, /* 0x382d */
            {8'h00}, /* 0x382c */
            {8'h00}, /* 0x382b */
            {8'h00}, /* 0x382a */
            {8'h00}, /* 0x3829 */
            {8'h00}, /* 0x3828 */
            {8'h00}, /* 0x3827 */
            {8'h00}, /* 0x3826 */
            {8'h00}, /* 0x3825 */
            {8'h00}, /* 0x3824 */
            {8'h00}, /* 0x3823 */
            {8'h00}, /* 0x3822 */
            {8'h00}, /* 0x3821 */
            {8'h00}, /* 0x3820 */
            {8'h00}, /* 0x381f */
            {8'h00}, /* 0x381e */
            {8'h00}, /* 0x381d */
            {8'h00}, /* 0x381c */
            {8'h00}, /* 0x381b */
            {8'h00}, /* 0x381a */
            {8'h00}, /* 0x3819 */
            {8'h00}, /* 0x3818 */
            {8'h00}, /* 0x3817 */
            {8'h00}, /* 0x3816 */
            {8'h00}, /* 0x3815 */
            {8'h00}, /* 0x3814 */
            {8'h00}, /* 0x3813 */
            {8'h00}, /* 0x3812 */
            {8'h00}, /* 0x3811 */
            {8'h00}, /* 0x3810 */
            {8'h00}, /* 0x380f */
            {8'h00}, /* 0x380e */
            {8'h00}, /* 0x380d */
            {8'h00}, /* 0x380c */
            {8'h00}, /* 0x380b */
            {8'h00}, /* 0x380a */
            {8'h00}, /* 0x3809 */
            {8'h00}, /* 0x3808 */
            {8'h00}, /* 0x3807 */
            {8'h00}, /* 0x3806 */
            {8'h00}, /* 0x3805 */
            {8'h00}, /* 0x3804 */
            {8'h00}, /* 0x3803 */
            {8'h00}, /* 0x3802 */
            {8'h00}, /* 0x3801 */
            {8'h00}, /* 0x3800 */
            {8'h00}, /* 0x37ff */
            {8'h00}, /* 0x37fe */
            {8'h00}, /* 0x37fd */
            {8'h00}, /* 0x37fc */
            {8'h00}, /* 0x37fb */
            {8'h00}, /* 0x37fa */
            {8'h00}, /* 0x37f9 */
            {8'h00}, /* 0x37f8 */
            {8'h00}, /* 0x37f7 */
            {8'h00}, /* 0x37f6 */
            {8'h00}, /* 0x37f5 */
            {8'h00}, /* 0x37f4 */
            {8'h00}, /* 0x37f3 */
            {8'h00}, /* 0x37f2 */
            {8'h00}, /* 0x37f1 */
            {8'h00}, /* 0x37f0 */
            {8'h00}, /* 0x37ef */
            {8'h00}, /* 0x37ee */
            {8'h00}, /* 0x37ed */
            {8'h00}, /* 0x37ec */
            {8'h00}, /* 0x37eb */
            {8'h00}, /* 0x37ea */
            {8'h00}, /* 0x37e9 */
            {8'h00}, /* 0x37e8 */
            {8'h00}, /* 0x37e7 */
            {8'h00}, /* 0x37e6 */
            {8'h00}, /* 0x37e5 */
            {8'h00}, /* 0x37e4 */
            {8'h00}, /* 0x37e3 */
            {8'h00}, /* 0x37e2 */
            {8'h00}, /* 0x37e1 */
            {8'h00}, /* 0x37e0 */
            {8'h00}, /* 0x37df */
            {8'h00}, /* 0x37de */
            {8'h00}, /* 0x37dd */
            {8'h00}, /* 0x37dc */
            {8'h00}, /* 0x37db */
            {8'h00}, /* 0x37da */
            {8'h00}, /* 0x37d9 */
            {8'h00}, /* 0x37d8 */
            {8'h00}, /* 0x37d7 */
            {8'h00}, /* 0x37d6 */
            {8'h00}, /* 0x37d5 */
            {8'h00}, /* 0x37d4 */
            {8'h00}, /* 0x37d3 */
            {8'h00}, /* 0x37d2 */
            {8'h00}, /* 0x37d1 */
            {8'h00}, /* 0x37d0 */
            {8'h00}, /* 0x37cf */
            {8'h00}, /* 0x37ce */
            {8'h00}, /* 0x37cd */
            {8'h00}, /* 0x37cc */
            {8'h00}, /* 0x37cb */
            {8'h00}, /* 0x37ca */
            {8'h00}, /* 0x37c9 */
            {8'h00}, /* 0x37c8 */
            {8'h00}, /* 0x37c7 */
            {8'h00}, /* 0x37c6 */
            {8'h00}, /* 0x37c5 */
            {8'h00}, /* 0x37c4 */
            {8'h00}, /* 0x37c3 */
            {8'h00}, /* 0x37c2 */
            {8'h00}, /* 0x37c1 */
            {8'h00}, /* 0x37c0 */
            {8'h00}, /* 0x37bf */
            {8'h00}, /* 0x37be */
            {8'h00}, /* 0x37bd */
            {8'h00}, /* 0x37bc */
            {8'h00}, /* 0x37bb */
            {8'h00}, /* 0x37ba */
            {8'h00}, /* 0x37b9 */
            {8'h00}, /* 0x37b8 */
            {8'h00}, /* 0x37b7 */
            {8'h00}, /* 0x37b6 */
            {8'h00}, /* 0x37b5 */
            {8'h00}, /* 0x37b4 */
            {8'h00}, /* 0x37b3 */
            {8'h00}, /* 0x37b2 */
            {8'h00}, /* 0x37b1 */
            {8'h00}, /* 0x37b0 */
            {8'h00}, /* 0x37af */
            {8'h00}, /* 0x37ae */
            {8'h00}, /* 0x37ad */
            {8'h00}, /* 0x37ac */
            {8'h00}, /* 0x37ab */
            {8'h00}, /* 0x37aa */
            {8'h00}, /* 0x37a9 */
            {8'h00}, /* 0x37a8 */
            {8'h00}, /* 0x37a7 */
            {8'h00}, /* 0x37a6 */
            {8'h00}, /* 0x37a5 */
            {8'h00}, /* 0x37a4 */
            {8'h00}, /* 0x37a3 */
            {8'h00}, /* 0x37a2 */
            {8'h00}, /* 0x37a1 */
            {8'h00}, /* 0x37a0 */
            {8'h00}, /* 0x379f */
            {8'h00}, /* 0x379e */
            {8'h00}, /* 0x379d */
            {8'h00}, /* 0x379c */
            {8'h00}, /* 0x379b */
            {8'h00}, /* 0x379a */
            {8'h00}, /* 0x3799 */
            {8'h00}, /* 0x3798 */
            {8'h00}, /* 0x3797 */
            {8'h00}, /* 0x3796 */
            {8'h00}, /* 0x3795 */
            {8'h00}, /* 0x3794 */
            {8'h00}, /* 0x3793 */
            {8'h00}, /* 0x3792 */
            {8'h00}, /* 0x3791 */
            {8'h00}, /* 0x3790 */
            {8'h00}, /* 0x378f */
            {8'h00}, /* 0x378e */
            {8'h00}, /* 0x378d */
            {8'h00}, /* 0x378c */
            {8'h00}, /* 0x378b */
            {8'h00}, /* 0x378a */
            {8'h00}, /* 0x3789 */
            {8'h00}, /* 0x3788 */
            {8'h00}, /* 0x3787 */
            {8'h00}, /* 0x3786 */
            {8'h00}, /* 0x3785 */
            {8'h00}, /* 0x3784 */
            {8'h00}, /* 0x3783 */
            {8'h00}, /* 0x3782 */
            {8'h00}, /* 0x3781 */
            {8'h00}, /* 0x3780 */
            {8'h00}, /* 0x377f */
            {8'h00}, /* 0x377e */
            {8'h00}, /* 0x377d */
            {8'h00}, /* 0x377c */
            {8'h00}, /* 0x377b */
            {8'h00}, /* 0x377a */
            {8'h00}, /* 0x3779 */
            {8'h00}, /* 0x3778 */
            {8'h00}, /* 0x3777 */
            {8'h00}, /* 0x3776 */
            {8'h00}, /* 0x3775 */
            {8'h00}, /* 0x3774 */
            {8'h00}, /* 0x3773 */
            {8'h00}, /* 0x3772 */
            {8'h00}, /* 0x3771 */
            {8'h00}, /* 0x3770 */
            {8'h00}, /* 0x376f */
            {8'h00}, /* 0x376e */
            {8'h00}, /* 0x376d */
            {8'h00}, /* 0x376c */
            {8'h00}, /* 0x376b */
            {8'h00}, /* 0x376a */
            {8'h00}, /* 0x3769 */
            {8'h00}, /* 0x3768 */
            {8'h00}, /* 0x3767 */
            {8'h00}, /* 0x3766 */
            {8'h00}, /* 0x3765 */
            {8'h00}, /* 0x3764 */
            {8'h00}, /* 0x3763 */
            {8'h00}, /* 0x3762 */
            {8'h00}, /* 0x3761 */
            {8'h00}, /* 0x3760 */
            {8'h00}, /* 0x375f */
            {8'h00}, /* 0x375e */
            {8'h00}, /* 0x375d */
            {8'h00}, /* 0x375c */
            {8'h00}, /* 0x375b */
            {8'h00}, /* 0x375a */
            {8'h00}, /* 0x3759 */
            {8'h00}, /* 0x3758 */
            {8'h00}, /* 0x3757 */
            {8'h00}, /* 0x3756 */
            {8'h00}, /* 0x3755 */
            {8'h00}, /* 0x3754 */
            {8'h00}, /* 0x3753 */
            {8'h00}, /* 0x3752 */
            {8'h00}, /* 0x3751 */
            {8'h00}, /* 0x3750 */
            {8'h00}, /* 0x374f */
            {8'h00}, /* 0x374e */
            {8'h00}, /* 0x374d */
            {8'h00}, /* 0x374c */
            {8'h00}, /* 0x374b */
            {8'h00}, /* 0x374a */
            {8'h00}, /* 0x3749 */
            {8'h00}, /* 0x3748 */
            {8'h00}, /* 0x3747 */
            {8'h00}, /* 0x3746 */
            {8'h00}, /* 0x3745 */
            {8'h00}, /* 0x3744 */
            {8'h00}, /* 0x3743 */
            {8'h00}, /* 0x3742 */
            {8'h00}, /* 0x3741 */
            {8'h00}, /* 0x3740 */
            {8'h00}, /* 0x373f */
            {8'h00}, /* 0x373e */
            {8'h00}, /* 0x373d */
            {8'h00}, /* 0x373c */
            {8'h00}, /* 0x373b */
            {8'h00}, /* 0x373a */
            {8'h00}, /* 0x3739 */
            {8'h00}, /* 0x3738 */
            {8'h00}, /* 0x3737 */
            {8'h00}, /* 0x3736 */
            {8'h00}, /* 0x3735 */
            {8'h00}, /* 0x3734 */
            {8'h00}, /* 0x3733 */
            {8'h00}, /* 0x3732 */
            {8'h00}, /* 0x3731 */
            {8'h00}, /* 0x3730 */
            {8'h00}, /* 0x372f */
            {8'h00}, /* 0x372e */
            {8'h00}, /* 0x372d */
            {8'h00}, /* 0x372c */
            {8'h00}, /* 0x372b */
            {8'h00}, /* 0x372a */
            {8'h00}, /* 0x3729 */
            {8'h00}, /* 0x3728 */
            {8'h00}, /* 0x3727 */
            {8'h00}, /* 0x3726 */
            {8'h00}, /* 0x3725 */
            {8'h00}, /* 0x3724 */
            {8'h00}, /* 0x3723 */
            {8'h00}, /* 0x3722 */
            {8'h00}, /* 0x3721 */
            {8'h00}, /* 0x3720 */
            {8'h00}, /* 0x371f */
            {8'h00}, /* 0x371e */
            {8'h00}, /* 0x371d */
            {8'h00}, /* 0x371c */
            {8'h00}, /* 0x371b */
            {8'h00}, /* 0x371a */
            {8'h00}, /* 0x3719 */
            {8'h00}, /* 0x3718 */
            {8'h00}, /* 0x3717 */
            {8'h00}, /* 0x3716 */
            {8'h00}, /* 0x3715 */
            {8'h00}, /* 0x3714 */
            {8'h00}, /* 0x3713 */
            {8'h00}, /* 0x3712 */
            {8'h00}, /* 0x3711 */
            {8'h00}, /* 0x3710 */
            {8'h00}, /* 0x370f */
            {8'h00}, /* 0x370e */
            {8'h00}, /* 0x370d */
            {8'h00}, /* 0x370c */
            {8'h00}, /* 0x370b */
            {8'h00}, /* 0x370a */
            {8'h00}, /* 0x3709 */
            {8'h00}, /* 0x3708 */
            {8'h00}, /* 0x3707 */
            {8'h00}, /* 0x3706 */
            {8'h00}, /* 0x3705 */
            {8'h00}, /* 0x3704 */
            {8'h00}, /* 0x3703 */
            {8'h00}, /* 0x3702 */
            {8'h00}, /* 0x3701 */
            {8'h00}, /* 0x3700 */
            {8'h00}, /* 0x36ff */
            {8'h00}, /* 0x36fe */
            {8'h00}, /* 0x36fd */
            {8'h00}, /* 0x36fc */
            {8'h00}, /* 0x36fb */
            {8'h00}, /* 0x36fa */
            {8'h00}, /* 0x36f9 */
            {8'h00}, /* 0x36f8 */
            {8'h00}, /* 0x36f7 */
            {8'h00}, /* 0x36f6 */
            {8'h00}, /* 0x36f5 */
            {8'h00}, /* 0x36f4 */
            {8'h00}, /* 0x36f3 */
            {8'h00}, /* 0x36f2 */
            {8'h00}, /* 0x36f1 */
            {8'h00}, /* 0x36f0 */
            {8'h00}, /* 0x36ef */
            {8'h00}, /* 0x36ee */
            {8'h00}, /* 0x36ed */
            {8'h00}, /* 0x36ec */
            {8'h00}, /* 0x36eb */
            {8'h00}, /* 0x36ea */
            {8'h00}, /* 0x36e9 */
            {8'h00}, /* 0x36e8 */
            {8'h00}, /* 0x36e7 */
            {8'h00}, /* 0x36e6 */
            {8'h00}, /* 0x36e5 */
            {8'h00}, /* 0x36e4 */
            {8'h00}, /* 0x36e3 */
            {8'h00}, /* 0x36e2 */
            {8'h00}, /* 0x36e1 */
            {8'h00}, /* 0x36e0 */
            {8'h00}, /* 0x36df */
            {8'h00}, /* 0x36de */
            {8'h00}, /* 0x36dd */
            {8'h00}, /* 0x36dc */
            {8'h00}, /* 0x36db */
            {8'h00}, /* 0x36da */
            {8'h00}, /* 0x36d9 */
            {8'h00}, /* 0x36d8 */
            {8'h00}, /* 0x36d7 */
            {8'h00}, /* 0x36d6 */
            {8'h00}, /* 0x36d5 */
            {8'h00}, /* 0x36d4 */
            {8'h00}, /* 0x36d3 */
            {8'h00}, /* 0x36d2 */
            {8'h00}, /* 0x36d1 */
            {8'h00}, /* 0x36d0 */
            {8'h00}, /* 0x36cf */
            {8'h00}, /* 0x36ce */
            {8'h00}, /* 0x36cd */
            {8'h00}, /* 0x36cc */
            {8'h00}, /* 0x36cb */
            {8'h00}, /* 0x36ca */
            {8'h00}, /* 0x36c9 */
            {8'h00}, /* 0x36c8 */
            {8'h00}, /* 0x36c7 */
            {8'h00}, /* 0x36c6 */
            {8'h00}, /* 0x36c5 */
            {8'h00}, /* 0x36c4 */
            {8'h00}, /* 0x36c3 */
            {8'h00}, /* 0x36c2 */
            {8'h00}, /* 0x36c1 */
            {8'h00}, /* 0x36c0 */
            {8'h00}, /* 0x36bf */
            {8'h00}, /* 0x36be */
            {8'h00}, /* 0x36bd */
            {8'h00}, /* 0x36bc */
            {8'h00}, /* 0x36bb */
            {8'h00}, /* 0x36ba */
            {8'h00}, /* 0x36b9 */
            {8'h00}, /* 0x36b8 */
            {8'h00}, /* 0x36b7 */
            {8'h00}, /* 0x36b6 */
            {8'h00}, /* 0x36b5 */
            {8'h00}, /* 0x36b4 */
            {8'h00}, /* 0x36b3 */
            {8'h00}, /* 0x36b2 */
            {8'h00}, /* 0x36b1 */
            {8'h00}, /* 0x36b0 */
            {8'h00}, /* 0x36af */
            {8'h00}, /* 0x36ae */
            {8'h00}, /* 0x36ad */
            {8'h00}, /* 0x36ac */
            {8'h00}, /* 0x36ab */
            {8'h00}, /* 0x36aa */
            {8'h00}, /* 0x36a9 */
            {8'h00}, /* 0x36a8 */
            {8'h00}, /* 0x36a7 */
            {8'h00}, /* 0x36a6 */
            {8'h00}, /* 0x36a5 */
            {8'h00}, /* 0x36a4 */
            {8'h00}, /* 0x36a3 */
            {8'h00}, /* 0x36a2 */
            {8'h00}, /* 0x36a1 */
            {8'h00}, /* 0x36a0 */
            {8'h00}, /* 0x369f */
            {8'h00}, /* 0x369e */
            {8'h00}, /* 0x369d */
            {8'h00}, /* 0x369c */
            {8'h00}, /* 0x369b */
            {8'h00}, /* 0x369a */
            {8'h00}, /* 0x3699 */
            {8'h00}, /* 0x3698 */
            {8'h00}, /* 0x3697 */
            {8'h00}, /* 0x3696 */
            {8'h00}, /* 0x3695 */
            {8'h00}, /* 0x3694 */
            {8'h00}, /* 0x3693 */
            {8'h00}, /* 0x3692 */
            {8'h00}, /* 0x3691 */
            {8'h00}, /* 0x3690 */
            {8'h00}, /* 0x368f */
            {8'h00}, /* 0x368e */
            {8'h00}, /* 0x368d */
            {8'h00}, /* 0x368c */
            {8'h00}, /* 0x368b */
            {8'h00}, /* 0x368a */
            {8'h00}, /* 0x3689 */
            {8'h00}, /* 0x3688 */
            {8'h00}, /* 0x3687 */
            {8'h00}, /* 0x3686 */
            {8'h00}, /* 0x3685 */
            {8'h00}, /* 0x3684 */
            {8'h00}, /* 0x3683 */
            {8'h00}, /* 0x3682 */
            {8'h00}, /* 0x3681 */
            {8'h00}, /* 0x3680 */
            {8'h00}, /* 0x367f */
            {8'h00}, /* 0x367e */
            {8'h00}, /* 0x367d */
            {8'h00}, /* 0x367c */
            {8'h00}, /* 0x367b */
            {8'h00}, /* 0x367a */
            {8'h00}, /* 0x3679 */
            {8'h00}, /* 0x3678 */
            {8'h00}, /* 0x3677 */
            {8'h00}, /* 0x3676 */
            {8'h00}, /* 0x3675 */
            {8'h00}, /* 0x3674 */
            {8'h00}, /* 0x3673 */
            {8'h00}, /* 0x3672 */
            {8'h00}, /* 0x3671 */
            {8'h00}, /* 0x3670 */
            {8'h00}, /* 0x366f */
            {8'h00}, /* 0x366e */
            {8'h00}, /* 0x366d */
            {8'h00}, /* 0x366c */
            {8'h00}, /* 0x366b */
            {8'h00}, /* 0x366a */
            {8'h00}, /* 0x3669 */
            {8'h00}, /* 0x3668 */
            {8'h00}, /* 0x3667 */
            {8'h00}, /* 0x3666 */
            {8'h00}, /* 0x3665 */
            {8'h00}, /* 0x3664 */
            {8'h00}, /* 0x3663 */
            {8'h00}, /* 0x3662 */
            {8'h00}, /* 0x3661 */
            {8'h00}, /* 0x3660 */
            {8'h00}, /* 0x365f */
            {8'h00}, /* 0x365e */
            {8'h00}, /* 0x365d */
            {8'h00}, /* 0x365c */
            {8'h00}, /* 0x365b */
            {8'h00}, /* 0x365a */
            {8'h00}, /* 0x3659 */
            {8'h00}, /* 0x3658 */
            {8'h00}, /* 0x3657 */
            {8'h00}, /* 0x3656 */
            {8'h00}, /* 0x3655 */
            {8'h00}, /* 0x3654 */
            {8'h00}, /* 0x3653 */
            {8'h00}, /* 0x3652 */
            {8'h00}, /* 0x3651 */
            {8'h00}, /* 0x3650 */
            {8'h00}, /* 0x364f */
            {8'h00}, /* 0x364e */
            {8'h00}, /* 0x364d */
            {8'h00}, /* 0x364c */
            {8'h00}, /* 0x364b */
            {8'h00}, /* 0x364a */
            {8'h00}, /* 0x3649 */
            {8'h00}, /* 0x3648 */
            {8'h00}, /* 0x3647 */
            {8'h00}, /* 0x3646 */
            {8'h00}, /* 0x3645 */
            {8'h00}, /* 0x3644 */
            {8'h00}, /* 0x3643 */
            {8'h00}, /* 0x3642 */
            {8'h00}, /* 0x3641 */
            {8'h00}, /* 0x3640 */
            {8'h00}, /* 0x363f */
            {8'h00}, /* 0x363e */
            {8'h00}, /* 0x363d */
            {8'h00}, /* 0x363c */
            {8'h00}, /* 0x363b */
            {8'h00}, /* 0x363a */
            {8'h00}, /* 0x3639 */
            {8'h00}, /* 0x3638 */
            {8'h00}, /* 0x3637 */
            {8'h00}, /* 0x3636 */
            {8'h00}, /* 0x3635 */
            {8'h00}, /* 0x3634 */
            {8'h00}, /* 0x3633 */
            {8'h00}, /* 0x3632 */
            {8'h00}, /* 0x3631 */
            {8'h00}, /* 0x3630 */
            {8'h00}, /* 0x362f */
            {8'h00}, /* 0x362e */
            {8'h00}, /* 0x362d */
            {8'h00}, /* 0x362c */
            {8'h00}, /* 0x362b */
            {8'h00}, /* 0x362a */
            {8'h00}, /* 0x3629 */
            {8'h00}, /* 0x3628 */
            {8'h00}, /* 0x3627 */
            {8'h00}, /* 0x3626 */
            {8'h00}, /* 0x3625 */
            {8'h00}, /* 0x3624 */
            {8'h00}, /* 0x3623 */
            {8'h00}, /* 0x3622 */
            {8'h00}, /* 0x3621 */
            {8'h00}, /* 0x3620 */
            {8'h00}, /* 0x361f */
            {8'h00}, /* 0x361e */
            {8'h00}, /* 0x361d */
            {8'h00}, /* 0x361c */
            {8'h00}, /* 0x361b */
            {8'h00}, /* 0x361a */
            {8'h00}, /* 0x3619 */
            {8'h00}, /* 0x3618 */
            {8'h00}, /* 0x3617 */
            {8'h00}, /* 0x3616 */
            {8'h00}, /* 0x3615 */
            {8'h00}, /* 0x3614 */
            {8'h00}, /* 0x3613 */
            {8'h00}, /* 0x3612 */
            {8'h00}, /* 0x3611 */
            {8'h00}, /* 0x3610 */
            {8'h00}, /* 0x360f */
            {8'h00}, /* 0x360e */
            {8'h00}, /* 0x360d */
            {8'h00}, /* 0x360c */
            {8'h00}, /* 0x360b */
            {8'h00}, /* 0x360a */
            {8'h00}, /* 0x3609 */
            {8'h00}, /* 0x3608 */
            {8'h00}, /* 0x3607 */
            {8'h00}, /* 0x3606 */
            {8'h00}, /* 0x3605 */
            {8'h00}, /* 0x3604 */
            {8'h00}, /* 0x3603 */
            {8'h00}, /* 0x3602 */
            {8'h00}, /* 0x3601 */
            {8'h00}, /* 0x3600 */
            {8'h00}, /* 0x35ff */
            {8'h00}, /* 0x35fe */
            {8'h00}, /* 0x35fd */
            {8'h00}, /* 0x35fc */
            {8'h00}, /* 0x35fb */
            {8'h00}, /* 0x35fa */
            {8'h00}, /* 0x35f9 */
            {8'h00}, /* 0x35f8 */
            {8'h00}, /* 0x35f7 */
            {8'h00}, /* 0x35f6 */
            {8'h00}, /* 0x35f5 */
            {8'h00}, /* 0x35f4 */
            {8'h00}, /* 0x35f3 */
            {8'h00}, /* 0x35f2 */
            {8'h00}, /* 0x35f1 */
            {8'h00}, /* 0x35f0 */
            {8'h00}, /* 0x35ef */
            {8'h00}, /* 0x35ee */
            {8'h00}, /* 0x35ed */
            {8'h00}, /* 0x35ec */
            {8'h00}, /* 0x35eb */
            {8'h00}, /* 0x35ea */
            {8'h00}, /* 0x35e9 */
            {8'h00}, /* 0x35e8 */
            {8'h00}, /* 0x35e7 */
            {8'h00}, /* 0x35e6 */
            {8'h00}, /* 0x35e5 */
            {8'h00}, /* 0x35e4 */
            {8'h00}, /* 0x35e3 */
            {8'h00}, /* 0x35e2 */
            {8'h00}, /* 0x35e1 */
            {8'h00}, /* 0x35e0 */
            {8'h00}, /* 0x35df */
            {8'h00}, /* 0x35de */
            {8'h00}, /* 0x35dd */
            {8'h00}, /* 0x35dc */
            {8'h00}, /* 0x35db */
            {8'h00}, /* 0x35da */
            {8'h00}, /* 0x35d9 */
            {8'h00}, /* 0x35d8 */
            {8'h00}, /* 0x35d7 */
            {8'h00}, /* 0x35d6 */
            {8'h00}, /* 0x35d5 */
            {8'h00}, /* 0x35d4 */
            {8'h00}, /* 0x35d3 */
            {8'h00}, /* 0x35d2 */
            {8'h00}, /* 0x35d1 */
            {8'h00}, /* 0x35d0 */
            {8'h00}, /* 0x35cf */
            {8'h00}, /* 0x35ce */
            {8'h00}, /* 0x35cd */
            {8'h00}, /* 0x35cc */
            {8'h00}, /* 0x35cb */
            {8'h00}, /* 0x35ca */
            {8'h00}, /* 0x35c9 */
            {8'h00}, /* 0x35c8 */
            {8'h00}, /* 0x35c7 */
            {8'h00}, /* 0x35c6 */
            {8'h00}, /* 0x35c5 */
            {8'h00}, /* 0x35c4 */
            {8'h00}, /* 0x35c3 */
            {8'h00}, /* 0x35c2 */
            {8'h00}, /* 0x35c1 */
            {8'h00}, /* 0x35c0 */
            {8'h00}, /* 0x35bf */
            {8'h00}, /* 0x35be */
            {8'h00}, /* 0x35bd */
            {8'h00}, /* 0x35bc */
            {8'h00}, /* 0x35bb */
            {8'h00}, /* 0x35ba */
            {8'h00}, /* 0x35b9 */
            {8'h00}, /* 0x35b8 */
            {8'h00}, /* 0x35b7 */
            {8'h00}, /* 0x35b6 */
            {8'h00}, /* 0x35b5 */
            {8'h00}, /* 0x35b4 */
            {8'h00}, /* 0x35b3 */
            {8'h00}, /* 0x35b2 */
            {8'h00}, /* 0x35b1 */
            {8'h00}, /* 0x35b0 */
            {8'h00}, /* 0x35af */
            {8'h00}, /* 0x35ae */
            {8'h00}, /* 0x35ad */
            {8'h00}, /* 0x35ac */
            {8'h00}, /* 0x35ab */
            {8'h00}, /* 0x35aa */
            {8'h00}, /* 0x35a9 */
            {8'h00}, /* 0x35a8 */
            {8'h00}, /* 0x35a7 */
            {8'h00}, /* 0x35a6 */
            {8'h00}, /* 0x35a5 */
            {8'h00}, /* 0x35a4 */
            {8'h00}, /* 0x35a3 */
            {8'h00}, /* 0x35a2 */
            {8'h00}, /* 0x35a1 */
            {8'h00}, /* 0x35a0 */
            {8'h00}, /* 0x359f */
            {8'h00}, /* 0x359e */
            {8'h00}, /* 0x359d */
            {8'h00}, /* 0x359c */
            {8'h00}, /* 0x359b */
            {8'h00}, /* 0x359a */
            {8'h00}, /* 0x3599 */
            {8'h00}, /* 0x3598 */
            {8'h00}, /* 0x3597 */
            {8'h00}, /* 0x3596 */
            {8'h00}, /* 0x3595 */
            {8'h00}, /* 0x3594 */
            {8'h00}, /* 0x3593 */
            {8'h00}, /* 0x3592 */
            {8'h00}, /* 0x3591 */
            {8'h00}, /* 0x3590 */
            {8'h00}, /* 0x358f */
            {8'h00}, /* 0x358e */
            {8'h00}, /* 0x358d */
            {8'h00}, /* 0x358c */
            {8'h00}, /* 0x358b */
            {8'h00}, /* 0x358a */
            {8'h00}, /* 0x3589 */
            {8'h00}, /* 0x3588 */
            {8'h00}, /* 0x3587 */
            {8'h00}, /* 0x3586 */
            {8'h00}, /* 0x3585 */
            {8'h00}, /* 0x3584 */
            {8'h00}, /* 0x3583 */
            {8'h00}, /* 0x3582 */
            {8'h00}, /* 0x3581 */
            {8'h00}, /* 0x3580 */
            {8'h00}, /* 0x357f */
            {8'h00}, /* 0x357e */
            {8'h00}, /* 0x357d */
            {8'h00}, /* 0x357c */
            {8'h00}, /* 0x357b */
            {8'h00}, /* 0x357a */
            {8'h00}, /* 0x3579 */
            {8'h00}, /* 0x3578 */
            {8'h00}, /* 0x3577 */
            {8'h00}, /* 0x3576 */
            {8'h00}, /* 0x3575 */
            {8'h00}, /* 0x3574 */
            {8'h00}, /* 0x3573 */
            {8'h00}, /* 0x3572 */
            {8'h00}, /* 0x3571 */
            {8'h00}, /* 0x3570 */
            {8'h00}, /* 0x356f */
            {8'h00}, /* 0x356e */
            {8'h00}, /* 0x356d */
            {8'h00}, /* 0x356c */
            {8'h00}, /* 0x356b */
            {8'h00}, /* 0x356a */
            {8'h00}, /* 0x3569 */
            {8'h00}, /* 0x3568 */
            {8'h00}, /* 0x3567 */
            {8'h00}, /* 0x3566 */
            {8'h00}, /* 0x3565 */
            {8'h00}, /* 0x3564 */
            {8'h00}, /* 0x3563 */
            {8'h00}, /* 0x3562 */
            {8'h00}, /* 0x3561 */
            {8'h00}, /* 0x3560 */
            {8'h00}, /* 0x355f */
            {8'h00}, /* 0x355e */
            {8'h00}, /* 0x355d */
            {8'h00}, /* 0x355c */
            {8'h00}, /* 0x355b */
            {8'h00}, /* 0x355a */
            {8'h00}, /* 0x3559 */
            {8'h00}, /* 0x3558 */
            {8'h00}, /* 0x3557 */
            {8'h00}, /* 0x3556 */
            {8'h00}, /* 0x3555 */
            {8'h00}, /* 0x3554 */
            {8'h00}, /* 0x3553 */
            {8'h00}, /* 0x3552 */
            {8'h00}, /* 0x3551 */
            {8'h00}, /* 0x3550 */
            {8'h00}, /* 0x354f */
            {8'h00}, /* 0x354e */
            {8'h00}, /* 0x354d */
            {8'h00}, /* 0x354c */
            {8'h00}, /* 0x354b */
            {8'h00}, /* 0x354a */
            {8'h00}, /* 0x3549 */
            {8'h00}, /* 0x3548 */
            {8'h00}, /* 0x3547 */
            {8'h00}, /* 0x3546 */
            {8'h00}, /* 0x3545 */
            {8'h00}, /* 0x3544 */
            {8'h00}, /* 0x3543 */
            {8'h00}, /* 0x3542 */
            {8'h00}, /* 0x3541 */
            {8'h00}, /* 0x3540 */
            {8'h00}, /* 0x353f */
            {8'h00}, /* 0x353e */
            {8'h00}, /* 0x353d */
            {8'h00}, /* 0x353c */
            {8'h00}, /* 0x353b */
            {8'h00}, /* 0x353a */
            {8'h00}, /* 0x3539 */
            {8'h00}, /* 0x3538 */
            {8'h00}, /* 0x3537 */
            {8'h00}, /* 0x3536 */
            {8'h00}, /* 0x3535 */
            {8'h00}, /* 0x3534 */
            {8'h00}, /* 0x3533 */
            {8'h00}, /* 0x3532 */
            {8'h00}, /* 0x3531 */
            {8'h00}, /* 0x3530 */
            {8'h00}, /* 0x352f */
            {8'h00}, /* 0x352e */
            {8'h00}, /* 0x352d */
            {8'h00}, /* 0x352c */
            {8'h00}, /* 0x352b */
            {8'h00}, /* 0x352a */
            {8'h00}, /* 0x3529 */
            {8'h00}, /* 0x3528 */
            {8'h00}, /* 0x3527 */
            {8'h00}, /* 0x3526 */
            {8'h00}, /* 0x3525 */
            {8'h00}, /* 0x3524 */
            {8'h00}, /* 0x3523 */
            {8'h00}, /* 0x3522 */
            {8'h00}, /* 0x3521 */
            {8'h00}, /* 0x3520 */
            {8'h00}, /* 0x351f */
            {8'h00}, /* 0x351e */
            {8'h00}, /* 0x351d */
            {8'h00}, /* 0x351c */
            {8'h00}, /* 0x351b */
            {8'h00}, /* 0x351a */
            {8'h00}, /* 0x3519 */
            {8'h00}, /* 0x3518 */
            {8'h00}, /* 0x3517 */
            {8'h00}, /* 0x3516 */
            {8'h00}, /* 0x3515 */
            {8'h00}, /* 0x3514 */
            {8'h00}, /* 0x3513 */
            {8'h00}, /* 0x3512 */
            {8'h00}, /* 0x3511 */
            {8'h00}, /* 0x3510 */
            {8'h00}, /* 0x350f */
            {8'h00}, /* 0x350e */
            {8'h00}, /* 0x350d */
            {8'h00}, /* 0x350c */
            {8'h00}, /* 0x350b */
            {8'h00}, /* 0x350a */
            {8'h00}, /* 0x3509 */
            {8'h00}, /* 0x3508 */
            {8'h00}, /* 0x3507 */
            {8'h00}, /* 0x3506 */
            {8'h00}, /* 0x3505 */
            {8'h00}, /* 0x3504 */
            {8'h00}, /* 0x3503 */
            {8'h00}, /* 0x3502 */
            {8'h00}, /* 0x3501 */
            {8'h00}, /* 0x3500 */
            {8'h00}, /* 0x34ff */
            {8'h00}, /* 0x34fe */
            {8'h00}, /* 0x34fd */
            {8'h00}, /* 0x34fc */
            {8'h00}, /* 0x34fb */
            {8'h00}, /* 0x34fa */
            {8'h00}, /* 0x34f9 */
            {8'h00}, /* 0x34f8 */
            {8'h00}, /* 0x34f7 */
            {8'h00}, /* 0x34f6 */
            {8'h00}, /* 0x34f5 */
            {8'h00}, /* 0x34f4 */
            {8'h00}, /* 0x34f3 */
            {8'h00}, /* 0x34f2 */
            {8'h00}, /* 0x34f1 */
            {8'h00}, /* 0x34f0 */
            {8'h00}, /* 0x34ef */
            {8'h00}, /* 0x34ee */
            {8'h00}, /* 0x34ed */
            {8'h00}, /* 0x34ec */
            {8'h00}, /* 0x34eb */
            {8'h00}, /* 0x34ea */
            {8'h00}, /* 0x34e9 */
            {8'h00}, /* 0x34e8 */
            {8'h00}, /* 0x34e7 */
            {8'h00}, /* 0x34e6 */
            {8'h00}, /* 0x34e5 */
            {8'h00}, /* 0x34e4 */
            {8'h00}, /* 0x34e3 */
            {8'h00}, /* 0x34e2 */
            {8'h00}, /* 0x34e1 */
            {8'h00}, /* 0x34e0 */
            {8'h00}, /* 0x34df */
            {8'h00}, /* 0x34de */
            {8'h00}, /* 0x34dd */
            {8'h00}, /* 0x34dc */
            {8'h00}, /* 0x34db */
            {8'h00}, /* 0x34da */
            {8'h00}, /* 0x34d9 */
            {8'h00}, /* 0x34d8 */
            {8'h00}, /* 0x34d7 */
            {8'h00}, /* 0x34d6 */
            {8'h00}, /* 0x34d5 */
            {8'h00}, /* 0x34d4 */
            {8'h00}, /* 0x34d3 */
            {8'h00}, /* 0x34d2 */
            {8'h00}, /* 0x34d1 */
            {8'h00}, /* 0x34d0 */
            {8'h00}, /* 0x34cf */
            {8'h00}, /* 0x34ce */
            {8'h00}, /* 0x34cd */
            {8'h00}, /* 0x34cc */
            {8'h00}, /* 0x34cb */
            {8'h00}, /* 0x34ca */
            {8'h00}, /* 0x34c9 */
            {8'h00}, /* 0x34c8 */
            {8'h00}, /* 0x34c7 */
            {8'h00}, /* 0x34c6 */
            {8'h00}, /* 0x34c5 */
            {8'h00}, /* 0x34c4 */
            {8'h00}, /* 0x34c3 */
            {8'h00}, /* 0x34c2 */
            {8'h00}, /* 0x34c1 */
            {8'h00}, /* 0x34c0 */
            {8'h00}, /* 0x34bf */
            {8'h00}, /* 0x34be */
            {8'h00}, /* 0x34bd */
            {8'h00}, /* 0x34bc */
            {8'h00}, /* 0x34bb */
            {8'h00}, /* 0x34ba */
            {8'h00}, /* 0x34b9 */
            {8'h00}, /* 0x34b8 */
            {8'h00}, /* 0x34b7 */
            {8'h00}, /* 0x34b6 */
            {8'h00}, /* 0x34b5 */
            {8'h00}, /* 0x34b4 */
            {8'h00}, /* 0x34b3 */
            {8'h00}, /* 0x34b2 */
            {8'h00}, /* 0x34b1 */
            {8'h00}, /* 0x34b0 */
            {8'h00}, /* 0x34af */
            {8'h00}, /* 0x34ae */
            {8'h00}, /* 0x34ad */
            {8'h00}, /* 0x34ac */
            {8'h00}, /* 0x34ab */
            {8'h00}, /* 0x34aa */
            {8'h00}, /* 0x34a9 */
            {8'h00}, /* 0x34a8 */
            {8'h00}, /* 0x34a7 */
            {8'h00}, /* 0x34a6 */
            {8'h00}, /* 0x34a5 */
            {8'h00}, /* 0x34a4 */
            {8'h00}, /* 0x34a3 */
            {8'h00}, /* 0x34a2 */
            {8'h00}, /* 0x34a1 */
            {8'h00}, /* 0x34a0 */
            {8'h00}, /* 0x349f */
            {8'h00}, /* 0x349e */
            {8'h00}, /* 0x349d */
            {8'h00}, /* 0x349c */
            {8'h00}, /* 0x349b */
            {8'h00}, /* 0x349a */
            {8'h00}, /* 0x3499 */
            {8'h00}, /* 0x3498 */
            {8'h00}, /* 0x3497 */
            {8'h00}, /* 0x3496 */
            {8'h00}, /* 0x3495 */
            {8'h00}, /* 0x3494 */
            {8'h00}, /* 0x3493 */
            {8'h00}, /* 0x3492 */
            {8'h00}, /* 0x3491 */
            {8'h00}, /* 0x3490 */
            {8'h00}, /* 0x348f */
            {8'h00}, /* 0x348e */
            {8'h00}, /* 0x348d */
            {8'h00}, /* 0x348c */
            {8'h00}, /* 0x348b */
            {8'h00}, /* 0x348a */
            {8'h00}, /* 0x3489 */
            {8'h00}, /* 0x3488 */
            {8'h00}, /* 0x3487 */
            {8'h00}, /* 0x3486 */
            {8'h00}, /* 0x3485 */
            {8'h00}, /* 0x3484 */
            {8'h00}, /* 0x3483 */
            {8'h00}, /* 0x3482 */
            {8'h00}, /* 0x3481 */
            {8'h00}, /* 0x3480 */
            {8'h00}, /* 0x347f */
            {8'h00}, /* 0x347e */
            {8'h00}, /* 0x347d */
            {8'h00}, /* 0x347c */
            {8'h00}, /* 0x347b */
            {8'h00}, /* 0x347a */
            {8'h00}, /* 0x3479 */
            {8'h00}, /* 0x3478 */
            {8'h00}, /* 0x3477 */
            {8'h00}, /* 0x3476 */
            {8'h00}, /* 0x3475 */
            {8'h00}, /* 0x3474 */
            {8'h00}, /* 0x3473 */
            {8'h00}, /* 0x3472 */
            {8'h00}, /* 0x3471 */
            {8'h00}, /* 0x3470 */
            {8'h00}, /* 0x346f */
            {8'h00}, /* 0x346e */
            {8'h00}, /* 0x346d */
            {8'h00}, /* 0x346c */
            {8'h00}, /* 0x346b */
            {8'h00}, /* 0x346a */
            {8'h00}, /* 0x3469 */
            {8'h00}, /* 0x3468 */
            {8'h00}, /* 0x3467 */
            {8'h00}, /* 0x3466 */
            {8'h00}, /* 0x3465 */
            {8'h00}, /* 0x3464 */
            {8'h00}, /* 0x3463 */
            {8'h00}, /* 0x3462 */
            {8'h00}, /* 0x3461 */
            {8'h00}, /* 0x3460 */
            {8'h00}, /* 0x345f */
            {8'h00}, /* 0x345e */
            {8'h00}, /* 0x345d */
            {8'h00}, /* 0x345c */
            {8'h00}, /* 0x345b */
            {8'h00}, /* 0x345a */
            {8'h00}, /* 0x3459 */
            {8'h00}, /* 0x3458 */
            {8'h00}, /* 0x3457 */
            {8'h00}, /* 0x3456 */
            {8'h00}, /* 0x3455 */
            {8'h00}, /* 0x3454 */
            {8'h00}, /* 0x3453 */
            {8'h00}, /* 0x3452 */
            {8'h00}, /* 0x3451 */
            {8'h00}, /* 0x3450 */
            {8'h00}, /* 0x344f */
            {8'h00}, /* 0x344e */
            {8'h00}, /* 0x344d */
            {8'h00}, /* 0x344c */
            {8'h00}, /* 0x344b */
            {8'h00}, /* 0x344a */
            {8'h00}, /* 0x3449 */
            {8'h00}, /* 0x3448 */
            {8'h00}, /* 0x3447 */
            {8'h00}, /* 0x3446 */
            {8'h00}, /* 0x3445 */
            {8'h00}, /* 0x3444 */
            {8'h00}, /* 0x3443 */
            {8'h00}, /* 0x3442 */
            {8'h00}, /* 0x3441 */
            {8'h00}, /* 0x3440 */
            {8'h00}, /* 0x343f */
            {8'h00}, /* 0x343e */
            {8'h00}, /* 0x343d */
            {8'h00}, /* 0x343c */
            {8'h00}, /* 0x343b */
            {8'h00}, /* 0x343a */
            {8'h00}, /* 0x3439 */
            {8'h00}, /* 0x3438 */
            {8'h00}, /* 0x3437 */
            {8'h00}, /* 0x3436 */
            {8'h00}, /* 0x3435 */
            {8'h00}, /* 0x3434 */
            {8'h00}, /* 0x3433 */
            {8'h00}, /* 0x3432 */
            {8'h00}, /* 0x3431 */
            {8'h00}, /* 0x3430 */
            {8'h00}, /* 0x342f */
            {8'h00}, /* 0x342e */
            {8'h00}, /* 0x342d */
            {8'h00}, /* 0x342c */
            {8'h00}, /* 0x342b */
            {8'h00}, /* 0x342a */
            {8'h00}, /* 0x3429 */
            {8'h00}, /* 0x3428 */
            {8'h00}, /* 0x3427 */
            {8'h00}, /* 0x3426 */
            {8'h00}, /* 0x3425 */
            {8'h00}, /* 0x3424 */
            {8'h00}, /* 0x3423 */
            {8'h00}, /* 0x3422 */
            {8'h00}, /* 0x3421 */
            {8'h00}, /* 0x3420 */
            {8'h00}, /* 0x341f */
            {8'h00}, /* 0x341e */
            {8'h00}, /* 0x341d */
            {8'h00}, /* 0x341c */
            {8'h00}, /* 0x341b */
            {8'h00}, /* 0x341a */
            {8'h00}, /* 0x3419 */
            {8'h00}, /* 0x3418 */
            {8'h00}, /* 0x3417 */
            {8'h00}, /* 0x3416 */
            {8'h00}, /* 0x3415 */
            {8'h00}, /* 0x3414 */
            {8'h00}, /* 0x3413 */
            {8'h00}, /* 0x3412 */
            {8'h00}, /* 0x3411 */
            {8'h00}, /* 0x3410 */
            {8'h00}, /* 0x340f */
            {8'h00}, /* 0x340e */
            {8'h00}, /* 0x340d */
            {8'h00}, /* 0x340c */
            {8'h00}, /* 0x340b */
            {8'h00}, /* 0x340a */
            {8'h00}, /* 0x3409 */
            {8'h00}, /* 0x3408 */
            {8'h00}, /* 0x3407 */
            {8'h00}, /* 0x3406 */
            {8'h00}, /* 0x3405 */
            {8'h00}, /* 0x3404 */
            {8'h00}, /* 0x3403 */
            {8'h00}, /* 0x3402 */
            {8'h00}, /* 0x3401 */
            {8'h00}, /* 0x3400 */
            {8'h00}, /* 0x33ff */
            {8'h00}, /* 0x33fe */
            {8'h00}, /* 0x33fd */
            {8'h00}, /* 0x33fc */
            {8'h00}, /* 0x33fb */
            {8'h00}, /* 0x33fa */
            {8'h00}, /* 0x33f9 */
            {8'h00}, /* 0x33f8 */
            {8'h00}, /* 0x33f7 */
            {8'h00}, /* 0x33f6 */
            {8'h00}, /* 0x33f5 */
            {8'h00}, /* 0x33f4 */
            {8'h00}, /* 0x33f3 */
            {8'h00}, /* 0x33f2 */
            {8'h00}, /* 0x33f1 */
            {8'h00}, /* 0x33f0 */
            {8'h00}, /* 0x33ef */
            {8'h00}, /* 0x33ee */
            {8'h00}, /* 0x33ed */
            {8'h00}, /* 0x33ec */
            {8'h00}, /* 0x33eb */
            {8'h00}, /* 0x33ea */
            {8'h00}, /* 0x33e9 */
            {8'h00}, /* 0x33e8 */
            {8'h00}, /* 0x33e7 */
            {8'h00}, /* 0x33e6 */
            {8'h00}, /* 0x33e5 */
            {8'h00}, /* 0x33e4 */
            {8'h00}, /* 0x33e3 */
            {8'h00}, /* 0x33e2 */
            {8'h00}, /* 0x33e1 */
            {8'h00}, /* 0x33e0 */
            {8'h00}, /* 0x33df */
            {8'h00}, /* 0x33de */
            {8'h00}, /* 0x33dd */
            {8'h00}, /* 0x33dc */
            {8'h00}, /* 0x33db */
            {8'h00}, /* 0x33da */
            {8'h00}, /* 0x33d9 */
            {8'h00}, /* 0x33d8 */
            {8'h00}, /* 0x33d7 */
            {8'h00}, /* 0x33d6 */
            {8'h00}, /* 0x33d5 */
            {8'h00}, /* 0x33d4 */
            {8'h00}, /* 0x33d3 */
            {8'h00}, /* 0x33d2 */
            {8'h00}, /* 0x33d1 */
            {8'h00}, /* 0x33d0 */
            {8'h00}, /* 0x33cf */
            {8'h00}, /* 0x33ce */
            {8'h00}, /* 0x33cd */
            {8'h00}, /* 0x33cc */
            {8'h00}, /* 0x33cb */
            {8'h00}, /* 0x33ca */
            {8'h00}, /* 0x33c9 */
            {8'h00}, /* 0x33c8 */
            {8'h00}, /* 0x33c7 */
            {8'h00}, /* 0x33c6 */
            {8'h00}, /* 0x33c5 */
            {8'h00}, /* 0x33c4 */
            {8'h00}, /* 0x33c3 */
            {8'h00}, /* 0x33c2 */
            {8'h00}, /* 0x33c1 */
            {8'h00}, /* 0x33c0 */
            {8'h00}, /* 0x33bf */
            {8'h00}, /* 0x33be */
            {8'h00}, /* 0x33bd */
            {8'h00}, /* 0x33bc */
            {8'h00}, /* 0x33bb */
            {8'h00}, /* 0x33ba */
            {8'h00}, /* 0x33b9 */
            {8'h00}, /* 0x33b8 */
            {8'h00}, /* 0x33b7 */
            {8'h00}, /* 0x33b6 */
            {8'h00}, /* 0x33b5 */
            {8'h00}, /* 0x33b4 */
            {8'h00}, /* 0x33b3 */
            {8'h00}, /* 0x33b2 */
            {8'h00}, /* 0x33b1 */
            {8'h00}, /* 0x33b0 */
            {8'h00}, /* 0x33af */
            {8'h00}, /* 0x33ae */
            {8'h00}, /* 0x33ad */
            {8'h00}, /* 0x33ac */
            {8'h00}, /* 0x33ab */
            {8'h00}, /* 0x33aa */
            {8'h00}, /* 0x33a9 */
            {8'h00}, /* 0x33a8 */
            {8'h00}, /* 0x33a7 */
            {8'h00}, /* 0x33a6 */
            {8'h00}, /* 0x33a5 */
            {8'h00}, /* 0x33a4 */
            {8'h00}, /* 0x33a3 */
            {8'h00}, /* 0x33a2 */
            {8'h00}, /* 0x33a1 */
            {8'h00}, /* 0x33a0 */
            {8'h00}, /* 0x339f */
            {8'h00}, /* 0x339e */
            {8'h00}, /* 0x339d */
            {8'h00}, /* 0x339c */
            {8'h00}, /* 0x339b */
            {8'h00}, /* 0x339a */
            {8'h00}, /* 0x3399 */
            {8'h00}, /* 0x3398 */
            {8'h00}, /* 0x3397 */
            {8'h00}, /* 0x3396 */
            {8'h00}, /* 0x3395 */
            {8'h00}, /* 0x3394 */
            {8'h00}, /* 0x3393 */
            {8'h00}, /* 0x3392 */
            {8'h00}, /* 0x3391 */
            {8'h00}, /* 0x3390 */
            {8'h00}, /* 0x338f */
            {8'h00}, /* 0x338e */
            {8'h00}, /* 0x338d */
            {8'h00}, /* 0x338c */
            {8'h00}, /* 0x338b */
            {8'h00}, /* 0x338a */
            {8'h00}, /* 0x3389 */
            {8'h00}, /* 0x3388 */
            {8'h00}, /* 0x3387 */
            {8'h00}, /* 0x3386 */
            {8'h00}, /* 0x3385 */
            {8'h00}, /* 0x3384 */
            {8'h00}, /* 0x3383 */
            {8'h00}, /* 0x3382 */
            {8'h00}, /* 0x3381 */
            {8'h00}, /* 0x3380 */
            {8'h00}, /* 0x337f */
            {8'h00}, /* 0x337e */
            {8'h00}, /* 0x337d */
            {8'h00}, /* 0x337c */
            {8'h00}, /* 0x337b */
            {8'h00}, /* 0x337a */
            {8'h00}, /* 0x3379 */
            {8'h00}, /* 0x3378 */
            {8'h00}, /* 0x3377 */
            {8'h00}, /* 0x3376 */
            {8'h00}, /* 0x3375 */
            {8'h00}, /* 0x3374 */
            {8'h00}, /* 0x3373 */
            {8'h00}, /* 0x3372 */
            {8'h00}, /* 0x3371 */
            {8'h00}, /* 0x3370 */
            {8'h00}, /* 0x336f */
            {8'h00}, /* 0x336e */
            {8'h00}, /* 0x336d */
            {8'h00}, /* 0x336c */
            {8'h00}, /* 0x336b */
            {8'h00}, /* 0x336a */
            {8'h00}, /* 0x3369 */
            {8'h00}, /* 0x3368 */
            {8'h00}, /* 0x3367 */
            {8'h00}, /* 0x3366 */
            {8'h00}, /* 0x3365 */
            {8'h00}, /* 0x3364 */
            {8'h00}, /* 0x3363 */
            {8'h00}, /* 0x3362 */
            {8'h00}, /* 0x3361 */
            {8'h00}, /* 0x3360 */
            {8'h00}, /* 0x335f */
            {8'h00}, /* 0x335e */
            {8'h00}, /* 0x335d */
            {8'h00}, /* 0x335c */
            {8'h00}, /* 0x335b */
            {8'h00}, /* 0x335a */
            {8'h00}, /* 0x3359 */
            {8'h00}, /* 0x3358 */
            {8'h00}, /* 0x3357 */
            {8'h00}, /* 0x3356 */
            {8'h00}, /* 0x3355 */
            {8'h00}, /* 0x3354 */
            {8'h00}, /* 0x3353 */
            {8'h00}, /* 0x3352 */
            {8'h00}, /* 0x3351 */
            {8'h00}, /* 0x3350 */
            {8'h00}, /* 0x334f */
            {8'h00}, /* 0x334e */
            {8'h00}, /* 0x334d */
            {8'h00}, /* 0x334c */
            {8'h00}, /* 0x334b */
            {8'h00}, /* 0x334a */
            {8'h00}, /* 0x3349 */
            {8'h00}, /* 0x3348 */
            {8'h00}, /* 0x3347 */
            {8'h00}, /* 0x3346 */
            {8'h00}, /* 0x3345 */
            {8'h00}, /* 0x3344 */
            {8'h00}, /* 0x3343 */
            {8'h00}, /* 0x3342 */
            {8'h00}, /* 0x3341 */
            {8'h00}, /* 0x3340 */
            {8'h00}, /* 0x333f */
            {8'h00}, /* 0x333e */
            {8'h00}, /* 0x333d */
            {8'h00}, /* 0x333c */
            {8'h00}, /* 0x333b */
            {8'h00}, /* 0x333a */
            {8'h00}, /* 0x3339 */
            {8'h00}, /* 0x3338 */
            {8'h00}, /* 0x3337 */
            {8'h00}, /* 0x3336 */
            {8'h00}, /* 0x3335 */
            {8'h00}, /* 0x3334 */
            {8'h00}, /* 0x3333 */
            {8'h00}, /* 0x3332 */
            {8'h00}, /* 0x3331 */
            {8'h00}, /* 0x3330 */
            {8'h00}, /* 0x332f */
            {8'h00}, /* 0x332e */
            {8'h00}, /* 0x332d */
            {8'h00}, /* 0x332c */
            {8'h00}, /* 0x332b */
            {8'h00}, /* 0x332a */
            {8'h00}, /* 0x3329 */
            {8'h00}, /* 0x3328 */
            {8'h00}, /* 0x3327 */
            {8'h00}, /* 0x3326 */
            {8'h00}, /* 0x3325 */
            {8'h00}, /* 0x3324 */
            {8'h00}, /* 0x3323 */
            {8'h00}, /* 0x3322 */
            {8'h00}, /* 0x3321 */
            {8'h00}, /* 0x3320 */
            {8'h00}, /* 0x331f */
            {8'h00}, /* 0x331e */
            {8'h00}, /* 0x331d */
            {8'h00}, /* 0x331c */
            {8'h00}, /* 0x331b */
            {8'h00}, /* 0x331a */
            {8'h00}, /* 0x3319 */
            {8'h00}, /* 0x3318 */
            {8'h00}, /* 0x3317 */
            {8'h00}, /* 0x3316 */
            {8'h00}, /* 0x3315 */
            {8'h00}, /* 0x3314 */
            {8'h00}, /* 0x3313 */
            {8'h00}, /* 0x3312 */
            {8'h00}, /* 0x3311 */
            {8'h00}, /* 0x3310 */
            {8'h00}, /* 0x330f */
            {8'h00}, /* 0x330e */
            {8'h00}, /* 0x330d */
            {8'h00}, /* 0x330c */
            {8'h00}, /* 0x330b */
            {8'h00}, /* 0x330a */
            {8'h00}, /* 0x3309 */
            {8'h00}, /* 0x3308 */
            {8'h00}, /* 0x3307 */
            {8'h00}, /* 0x3306 */
            {8'h00}, /* 0x3305 */
            {8'h00}, /* 0x3304 */
            {8'h00}, /* 0x3303 */
            {8'h00}, /* 0x3302 */
            {8'h00}, /* 0x3301 */
            {8'h00}, /* 0x3300 */
            {8'h00}, /* 0x32ff */
            {8'h00}, /* 0x32fe */
            {8'h00}, /* 0x32fd */
            {8'h00}, /* 0x32fc */
            {8'h00}, /* 0x32fb */
            {8'h00}, /* 0x32fa */
            {8'h00}, /* 0x32f9 */
            {8'h00}, /* 0x32f8 */
            {8'h00}, /* 0x32f7 */
            {8'h00}, /* 0x32f6 */
            {8'h00}, /* 0x32f5 */
            {8'h00}, /* 0x32f4 */
            {8'h00}, /* 0x32f3 */
            {8'h00}, /* 0x32f2 */
            {8'h00}, /* 0x32f1 */
            {8'h00}, /* 0x32f0 */
            {8'h00}, /* 0x32ef */
            {8'h00}, /* 0x32ee */
            {8'h00}, /* 0x32ed */
            {8'h00}, /* 0x32ec */
            {8'h00}, /* 0x32eb */
            {8'h00}, /* 0x32ea */
            {8'h00}, /* 0x32e9 */
            {8'h00}, /* 0x32e8 */
            {8'h00}, /* 0x32e7 */
            {8'h00}, /* 0x32e6 */
            {8'h00}, /* 0x32e5 */
            {8'h00}, /* 0x32e4 */
            {8'h00}, /* 0x32e3 */
            {8'h00}, /* 0x32e2 */
            {8'h00}, /* 0x32e1 */
            {8'h00}, /* 0x32e0 */
            {8'h00}, /* 0x32df */
            {8'h00}, /* 0x32de */
            {8'h00}, /* 0x32dd */
            {8'h00}, /* 0x32dc */
            {8'h00}, /* 0x32db */
            {8'h00}, /* 0x32da */
            {8'h00}, /* 0x32d9 */
            {8'h00}, /* 0x32d8 */
            {8'h00}, /* 0x32d7 */
            {8'h00}, /* 0x32d6 */
            {8'h00}, /* 0x32d5 */
            {8'h00}, /* 0x32d4 */
            {8'h00}, /* 0x32d3 */
            {8'h00}, /* 0x32d2 */
            {8'h00}, /* 0x32d1 */
            {8'h00}, /* 0x32d0 */
            {8'h00}, /* 0x32cf */
            {8'h00}, /* 0x32ce */
            {8'h00}, /* 0x32cd */
            {8'h00}, /* 0x32cc */
            {8'h00}, /* 0x32cb */
            {8'h00}, /* 0x32ca */
            {8'h00}, /* 0x32c9 */
            {8'h00}, /* 0x32c8 */
            {8'h00}, /* 0x32c7 */
            {8'h00}, /* 0x32c6 */
            {8'h00}, /* 0x32c5 */
            {8'h00}, /* 0x32c4 */
            {8'h00}, /* 0x32c3 */
            {8'h00}, /* 0x32c2 */
            {8'h00}, /* 0x32c1 */
            {8'h00}, /* 0x32c0 */
            {8'h00}, /* 0x32bf */
            {8'h00}, /* 0x32be */
            {8'h00}, /* 0x32bd */
            {8'h00}, /* 0x32bc */
            {8'h00}, /* 0x32bb */
            {8'h00}, /* 0x32ba */
            {8'h00}, /* 0x32b9 */
            {8'h00}, /* 0x32b8 */
            {8'h00}, /* 0x32b7 */
            {8'h00}, /* 0x32b6 */
            {8'h00}, /* 0x32b5 */
            {8'h00}, /* 0x32b4 */
            {8'h00}, /* 0x32b3 */
            {8'h00}, /* 0x32b2 */
            {8'h00}, /* 0x32b1 */
            {8'h00}, /* 0x32b0 */
            {8'h00}, /* 0x32af */
            {8'h00}, /* 0x32ae */
            {8'h00}, /* 0x32ad */
            {8'h00}, /* 0x32ac */
            {8'h00}, /* 0x32ab */
            {8'h00}, /* 0x32aa */
            {8'h00}, /* 0x32a9 */
            {8'h00}, /* 0x32a8 */
            {8'h00}, /* 0x32a7 */
            {8'h00}, /* 0x32a6 */
            {8'h00}, /* 0x32a5 */
            {8'h00}, /* 0x32a4 */
            {8'h00}, /* 0x32a3 */
            {8'h00}, /* 0x32a2 */
            {8'h00}, /* 0x32a1 */
            {8'h00}, /* 0x32a0 */
            {8'h00}, /* 0x329f */
            {8'h00}, /* 0x329e */
            {8'h00}, /* 0x329d */
            {8'h00}, /* 0x329c */
            {8'h00}, /* 0x329b */
            {8'h00}, /* 0x329a */
            {8'h00}, /* 0x3299 */
            {8'h00}, /* 0x3298 */
            {8'h00}, /* 0x3297 */
            {8'h00}, /* 0x3296 */
            {8'h00}, /* 0x3295 */
            {8'h00}, /* 0x3294 */
            {8'h00}, /* 0x3293 */
            {8'h00}, /* 0x3292 */
            {8'h00}, /* 0x3291 */
            {8'h00}, /* 0x3290 */
            {8'h00}, /* 0x328f */
            {8'h00}, /* 0x328e */
            {8'h00}, /* 0x328d */
            {8'h00}, /* 0x328c */
            {8'h00}, /* 0x328b */
            {8'h00}, /* 0x328a */
            {8'h00}, /* 0x3289 */
            {8'h00}, /* 0x3288 */
            {8'h00}, /* 0x3287 */
            {8'h00}, /* 0x3286 */
            {8'h00}, /* 0x3285 */
            {8'h00}, /* 0x3284 */
            {8'h00}, /* 0x3283 */
            {8'h00}, /* 0x3282 */
            {8'h00}, /* 0x3281 */
            {8'h00}, /* 0x3280 */
            {8'h00}, /* 0x327f */
            {8'h00}, /* 0x327e */
            {8'h00}, /* 0x327d */
            {8'h00}, /* 0x327c */
            {8'h00}, /* 0x327b */
            {8'h00}, /* 0x327a */
            {8'h00}, /* 0x3279 */
            {8'h00}, /* 0x3278 */
            {8'h00}, /* 0x3277 */
            {8'h00}, /* 0x3276 */
            {8'h00}, /* 0x3275 */
            {8'h00}, /* 0x3274 */
            {8'h00}, /* 0x3273 */
            {8'h00}, /* 0x3272 */
            {8'h00}, /* 0x3271 */
            {8'h00}, /* 0x3270 */
            {8'h00}, /* 0x326f */
            {8'h00}, /* 0x326e */
            {8'h00}, /* 0x326d */
            {8'h00}, /* 0x326c */
            {8'h00}, /* 0x326b */
            {8'h00}, /* 0x326a */
            {8'h00}, /* 0x3269 */
            {8'h00}, /* 0x3268 */
            {8'h00}, /* 0x3267 */
            {8'h00}, /* 0x3266 */
            {8'h00}, /* 0x3265 */
            {8'h00}, /* 0x3264 */
            {8'h00}, /* 0x3263 */
            {8'h00}, /* 0x3262 */
            {8'h00}, /* 0x3261 */
            {8'h00}, /* 0x3260 */
            {8'h00}, /* 0x325f */
            {8'h00}, /* 0x325e */
            {8'h00}, /* 0x325d */
            {8'h00}, /* 0x325c */
            {8'h00}, /* 0x325b */
            {8'h00}, /* 0x325a */
            {8'h00}, /* 0x3259 */
            {8'h00}, /* 0x3258 */
            {8'h00}, /* 0x3257 */
            {8'h00}, /* 0x3256 */
            {8'h00}, /* 0x3255 */
            {8'h00}, /* 0x3254 */
            {8'h00}, /* 0x3253 */
            {8'h00}, /* 0x3252 */
            {8'h00}, /* 0x3251 */
            {8'h00}, /* 0x3250 */
            {8'h00}, /* 0x324f */
            {8'h00}, /* 0x324e */
            {8'h00}, /* 0x324d */
            {8'h00}, /* 0x324c */
            {8'h00}, /* 0x324b */
            {8'h00}, /* 0x324a */
            {8'h00}, /* 0x3249 */
            {8'h00}, /* 0x3248 */
            {8'h00}, /* 0x3247 */
            {8'h00}, /* 0x3246 */
            {8'h00}, /* 0x3245 */
            {8'h00}, /* 0x3244 */
            {8'h00}, /* 0x3243 */
            {8'h00}, /* 0x3242 */
            {8'h00}, /* 0x3241 */
            {8'h00}, /* 0x3240 */
            {8'h00}, /* 0x323f */
            {8'h00}, /* 0x323e */
            {8'h00}, /* 0x323d */
            {8'h00}, /* 0x323c */
            {8'h00}, /* 0x323b */
            {8'h00}, /* 0x323a */
            {8'h00}, /* 0x3239 */
            {8'h00}, /* 0x3238 */
            {8'h00}, /* 0x3237 */
            {8'h00}, /* 0x3236 */
            {8'h00}, /* 0x3235 */
            {8'h00}, /* 0x3234 */
            {8'h00}, /* 0x3233 */
            {8'h00}, /* 0x3232 */
            {8'h00}, /* 0x3231 */
            {8'h00}, /* 0x3230 */
            {8'h00}, /* 0x322f */
            {8'h00}, /* 0x322e */
            {8'h00}, /* 0x322d */
            {8'h00}, /* 0x322c */
            {8'h00}, /* 0x322b */
            {8'h00}, /* 0x322a */
            {8'h00}, /* 0x3229 */
            {8'h00}, /* 0x3228 */
            {8'h00}, /* 0x3227 */
            {8'h00}, /* 0x3226 */
            {8'h00}, /* 0x3225 */
            {8'h00}, /* 0x3224 */
            {8'h00}, /* 0x3223 */
            {8'h00}, /* 0x3222 */
            {8'h00}, /* 0x3221 */
            {8'h00}, /* 0x3220 */
            {8'h00}, /* 0x321f */
            {8'h00}, /* 0x321e */
            {8'h00}, /* 0x321d */
            {8'h00}, /* 0x321c */
            {8'h00}, /* 0x321b */
            {8'h00}, /* 0x321a */
            {8'h00}, /* 0x3219 */
            {8'h00}, /* 0x3218 */
            {8'h00}, /* 0x3217 */
            {8'h00}, /* 0x3216 */
            {8'h00}, /* 0x3215 */
            {8'h00}, /* 0x3214 */
            {8'h00}, /* 0x3213 */
            {8'h00}, /* 0x3212 */
            {8'h00}, /* 0x3211 */
            {8'h00}, /* 0x3210 */
            {8'h00}, /* 0x320f */
            {8'h00}, /* 0x320e */
            {8'h00}, /* 0x320d */
            {8'h00}, /* 0x320c */
            {8'h00}, /* 0x320b */
            {8'h00}, /* 0x320a */
            {8'h00}, /* 0x3209 */
            {8'h00}, /* 0x3208 */
            {8'h00}, /* 0x3207 */
            {8'h00}, /* 0x3206 */
            {8'h00}, /* 0x3205 */
            {8'h00}, /* 0x3204 */
            {8'h00}, /* 0x3203 */
            {8'h00}, /* 0x3202 */
            {8'h00}, /* 0x3201 */
            {8'h00}, /* 0x3200 */
            {8'h00}, /* 0x31ff */
            {8'h00}, /* 0x31fe */
            {8'h00}, /* 0x31fd */
            {8'h00}, /* 0x31fc */
            {8'h00}, /* 0x31fb */
            {8'h00}, /* 0x31fa */
            {8'h00}, /* 0x31f9 */
            {8'h00}, /* 0x31f8 */
            {8'h00}, /* 0x31f7 */
            {8'h00}, /* 0x31f6 */
            {8'h00}, /* 0x31f5 */
            {8'h00}, /* 0x31f4 */
            {8'h00}, /* 0x31f3 */
            {8'h00}, /* 0x31f2 */
            {8'h00}, /* 0x31f1 */
            {8'h00}, /* 0x31f0 */
            {8'h00}, /* 0x31ef */
            {8'h00}, /* 0x31ee */
            {8'h00}, /* 0x31ed */
            {8'h00}, /* 0x31ec */
            {8'h00}, /* 0x31eb */
            {8'h00}, /* 0x31ea */
            {8'h00}, /* 0x31e9 */
            {8'h00}, /* 0x31e8 */
            {8'h00}, /* 0x31e7 */
            {8'h00}, /* 0x31e6 */
            {8'h00}, /* 0x31e5 */
            {8'h00}, /* 0x31e4 */
            {8'h00}, /* 0x31e3 */
            {8'h00}, /* 0x31e2 */
            {8'h00}, /* 0x31e1 */
            {8'h00}, /* 0x31e0 */
            {8'h00}, /* 0x31df */
            {8'h00}, /* 0x31de */
            {8'h00}, /* 0x31dd */
            {8'h00}, /* 0x31dc */
            {8'h00}, /* 0x31db */
            {8'h00}, /* 0x31da */
            {8'h00}, /* 0x31d9 */
            {8'h00}, /* 0x31d8 */
            {8'h00}, /* 0x31d7 */
            {8'h00}, /* 0x31d6 */
            {8'h00}, /* 0x31d5 */
            {8'h00}, /* 0x31d4 */
            {8'h00}, /* 0x31d3 */
            {8'h00}, /* 0x31d2 */
            {8'h00}, /* 0x31d1 */
            {8'h00}, /* 0x31d0 */
            {8'h00}, /* 0x31cf */
            {8'h00}, /* 0x31ce */
            {8'h00}, /* 0x31cd */
            {8'h00}, /* 0x31cc */
            {8'h00}, /* 0x31cb */
            {8'h00}, /* 0x31ca */
            {8'h00}, /* 0x31c9 */
            {8'h00}, /* 0x31c8 */
            {8'h00}, /* 0x31c7 */
            {8'h00}, /* 0x31c6 */
            {8'h00}, /* 0x31c5 */
            {8'h00}, /* 0x31c4 */
            {8'h00}, /* 0x31c3 */
            {8'h00}, /* 0x31c2 */
            {8'h00}, /* 0x31c1 */
            {8'h00}, /* 0x31c0 */
            {8'h00}, /* 0x31bf */
            {8'h00}, /* 0x31be */
            {8'h00}, /* 0x31bd */
            {8'h00}, /* 0x31bc */
            {8'h00}, /* 0x31bb */
            {8'h00}, /* 0x31ba */
            {8'h00}, /* 0x31b9 */
            {8'h00}, /* 0x31b8 */
            {8'h00}, /* 0x31b7 */
            {8'h00}, /* 0x31b6 */
            {8'h00}, /* 0x31b5 */
            {8'h00}, /* 0x31b4 */
            {8'h00}, /* 0x31b3 */
            {8'h00}, /* 0x31b2 */
            {8'h00}, /* 0x31b1 */
            {8'h00}, /* 0x31b0 */
            {8'h00}, /* 0x31af */
            {8'h00}, /* 0x31ae */
            {8'h00}, /* 0x31ad */
            {8'h00}, /* 0x31ac */
            {8'h00}, /* 0x31ab */
            {8'h00}, /* 0x31aa */
            {8'h00}, /* 0x31a9 */
            {8'h00}, /* 0x31a8 */
            {8'h00}, /* 0x31a7 */
            {8'h00}, /* 0x31a6 */
            {8'h00}, /* 0x31a5 */
            {8'h00}, /* 0x31a4 */
            {8'h00}, /* 0x31a3 */
            {8'h00}, /* 0x31a2 */
            {8'h00}, /* 0x31a1 */
            {8'h00}, /* 0x31a0 */
            {8'h00}, /* 0x319f */
            {8'h00}, /* 0x319e */
            {8'h00}, /* 0x319d */
            {8'h00}, /* 0x319c */
            {8'h00}, /* 0x319b */
            {8'h00}, /* 0x319a */
            {8'h00}, /* 0x3199 */
            {8'h00}, /* 0x3198 */
            {8'h00}, /* 0x3197 */
            {8'h00}, /* 0x3196 */
            {8'h00}, /* 0x3195 */
            {8'h00}, /* 0x3194 */
            {8'h00}, /* 0x3193 */
            {8'h00}, /* 0x3192 */
            {8'h00}, /* 0x3191 */
            {8'h00}, /* 0x3190 */
            {8'h00}, /* 0x318f */
            {8'h00}, /* 0x318e */
            {8'h00}, /* 0x318d */
            {8'h00}, /* 0x318c */
            {8'h00}, /* 0x318b */
            {8'h00}, /* 0x318a */
            {8'h00}, /* 0x3189 */
            {8'h00}, /* 0x3188 */
            {8'h00}, /* 0x3187 */
            {8'h00}, /* 0x3186 */
            {8'h00}, /* 0x3185 */
            {8'h00}, /* 0x3184 */
            {8'h00}, /* 0x3183 */
            {8'h00}, /* 0x3182 */
            {8'h00}, /* 0x3181 */
            {8'h00}, /* 0x3180 */
            {8'h00}, /* 0x317f */
            {8'h00}, /* 0x317e */
            {8'h00}, /* 0x317d */
            {8'h00}, /* 0x317c */
            {8'h00}, /* 0x317b */
            {8'h00}, /* 0x317a */
            {8'h00}, /* 0x3179 */
            {8'h00}, /* 0x3178 */
            {8'h00}, /* 0x3177 */
            {8'h00}, /* 0x3176 */
            {8'h00}, /* 0x3175 */
            {8'h00}, /* 0x3174 */
            {8'h00}, /* 0x3173 */
            {8'h00}, /* 0x3172 */
            {8'h00}, /* 0x3171 */
            {8'h00}, /* 0x3170 */
            {8'h00}, /* 0x316f */
            {8'h00}, /* 0x316e */
            {8'h00}, /* 0x316d */
            {8'h00}, /* 0x316c */
            {8'h00}, /* 0x316b */
            {8'h00}, /* 0x316a */
            {8'h00}, /* 0x3169 */
            {8'h00}, /* 0x3168 */
            {8'h00}, /* 0x3167 */
            {8'h00}, /* 0x3166 */
            {8'h00}, /* 0x3165 */
            {8'h00}, /* 0x3164 */
            {8'h00}, /* 0x3163 */
            {8'h00}, /* 0x3162 */
            {8'h00}, /* 0x3161 */
            {8'h00}, /* 0x3160 */
            {8'h00}, /* 0x315f */
            {8'h00}, /* 0x315e */
            {8'h00}, /* 0x315d */
            {8'h00}, /* 0x315c */
            {8'h00}, /* 0x315b */
            {8'h00}, /* 0x315a */
            {8'h00}, /* 0x3159 */
            {8'h00}, /* 0x3158 */
            {8'h00}, /* 0x3157 */
            {8'h00}, /* 0x3156 */
            {8'h00}, /* 0x3155 */
            {8'h00}, /* 0x3154 */
            {8'h00}, /* 0x3153 */
            {8'h00}, /* 0x3152 */
            {8'h00}, /* 0x3151 */
            {8'h00}, /* 0x3150 */
            {8'h00}, /* 0x314f */
            {8'h00}, /* 0x314e */
            {8'h00}, /* 0x314d */
            {8'h00}, /* 0x314c */
            {8'h00}, /* 0x314b */
            {8'h00}, /* 0x314a */
            {8'h00}, /* 0x3149 */
            {8'h00}, /* 0x3148 */
            {8'h00}, /* 0x3147 */
            {8'h00}, /* 0x3146 */
            {8'h00}, /* 0x3145 */
            {8'h00}, /* 0x3144 */
            {8'h00}, /* 0x3143 */
            {8'h00}, /* 0x3142 */
            {8'h00}, /* 0x3141 */
            {8'h00}, /* 0x3140 */
            {8'h00}, /* 0x313f */
            {8'h00}, /* 0x313e */
            {8'h00}, /* 0x313d */
            {8'h00}, /* 0x313c */
            {8'h00}, /* 0x313b */
            {8'h00}, /* 0x313a */
            {8'h00}, /* 0x3139 */
            {8'h00}, /* 0x3138 */
            {8'h00}, /* 0x3137 */
            {8'h00}, /* 0x3136 */
            {8'h00}, /* 0x3135 */
            {8'h00}, /* 0x3134 */
            {8'h00}, /* 0x3133 */
            {8'h00}, /* 0x3132 */
            {8'h00}, /* 0x3131 */
            {8'h00}, /* 0x3130 */
            {8'h00}, /* 0x312f */
            {8'h00}, /* 0x312e */
            {8'h00}, /* 0x312d */
            {8'h00}, /* 0x312c */
            {8'h00}, /* 0x312b */
            {8'h00}, /* 0x312a */
            {8'h00}, /* 0x3129 */
            {8'h00}, /* 0x3128 */
            {8'h00}, /* 0x3127 */
            {8'h00}, /* 0x3126 */
            {8'h00}, /* 0x3125 */
            {8'h00}, /* 0x3124 */
            {8'h00}, /* 0x3123 */
            {8'h00}, /* 0x3122 */
            {8'h00}, /* 0x3121 */
            {8'h00}, /* 0x3120 */
            {8'h00}, /* 0x311f */
            {8'h00}, /* 0x311e */
            {8'h00}, /* 0x311d */
            {8'h00}, /* 0x311c */
            {8'h00}, /* 0x311b */
            {8'h00}, /* 0x311a */
            {8'h00}, /* 0x3119 */
            {8'h00}, /* 0x3118 */
            {8'h00}, /* 0x3117 */
            {8'h00}, /* 0x3116 */
            {8'h00}, /* 0x3115 */
            {8'h00}, /* 0x3114 */
            {8'h00}, /* 0x3113 */
            {8'h00}, /* 0x3112 */
            {8'h00}, /* 0x3111 */
            {8'h00}, /* 0x3110 */
            {8'h00}, /* 0x310f */
            {8'h00}, /* 0x310e */
            {8'h00}, /* 0x310d */
            {8'h00}, /* 0x310c */
            {8'h00}, /* 0x310b */
            {8'h00}, /* 0x310a */
            {8'h00}, /* 0x3109 */
            {8'h00}, /* 0x3108 */
            {8'h00}, /* 0x3107 */
            {8'h00}, /* 0x3106 */
            {8'h00}, /* 0x3105 */
            {8'h00}, /* 0x3104 */
            {8'h00}, /* 0x3103 */
            {8'h00}, /* 0x3102 */
            {8'h00}, /* 0x3101 */
            {8'h00}, /* 0x3100 */
            {8'h00}, /* 0x30ff */
            {8'h00}, /* 0x30fe */
            {8'h00}, /* 0x30fd */
            {8'h00}, /* 0x30fc */
            {8'h00}, /* 0x30fb */
            {8'h00}, /* 0x30fa */
            {8'h00}, /* 0x30f9 */
            {8'h00}, /* 0x30f8 */
            {8'h00}, /* 0x30f7 */
            {8'h00}, /* 0x30f6 */
            {8'h00}, /* 0x30f5 */
            {8'h00}, /* 0x30f4 */
            {8'h00}, /* 0x30f3 */
            {8'h00}, /* 0x30f2 */
            {8'h00}, /* 0x30f1 */
            {8'h00}, /* 0x30f0 */
            {8'h00}, /* 0x30ef */
            {8'h00}, /* 0x30ee */
            {8'h00}, /* 0x30ed */
            {8'h00}, /* 0x30ec */
            {8'h00}, /* 0x30eb */
            {8'h00}, /* 0x30ea */
            {8'h00}, /* 0x30e9 */
            {8'h00}, /* 0x30e8 */
            {8'h00}, /* 0x30e7 */
            {8'h00}, /* 0x30e6 */
            {8'h00}, /* 0x30e5 */
            {8'h00}, /* 0x30e4 */
            {8'h00}, /* 0x30e3 */
            {8'h00}, /* 0x30e2 */
            {8'h00}, /* 0x30e1 */
            {8'h00}, /* 0x30e0 */
            {8'h00}, /* 0x30df */
            {8'h00}, /* 0x30de */
            {8'h00}, /* 0x30dd */
            {8'h00}, /* 0x30dc */
            {8'h00}, /* 0x30db */
            {8'h00}, /* 0x30da */
            {8'h00}, /* 0x30d9 */
            {8'h00}, /* 0x30d8 */
            {8'h00}, /* 0x30d7 */
            {8'h00}, /* 0x30d6 */
            {8'h00}, /* 0x30d5 */
            {8'h00}, /* 0x30d4 */
            {8'h00}, /* 0x30d3 */
            {8'h00}, /* 0x30d2 */
            {8'h00}, /* 0x30d1 */
            {8'h00}, /* 0x30d0 */
            {8'h00}, /* 0x30cf */
            {8'h00}, /* 0x30ce */
            {8'h00}, /* 0x30cd */
            {8'h00}, /* 0x30cc */
            {8'h00}, /* 0x30cb */
            {8'h00}, /* 0x30ca */
            {8'h00}, /* 0x30c9 */
            {8'h00}, /* 0x30c8 */
            {8'h00}, /* 0x30c7 */
            {8'h00}, /* 0x30c6 */
            {8'h00}, /* 0x30c5 */
            {8'h00}, /* 0x30c4 */
            {8'h00}, /* 0x30c3 */
            {8'h00}, /* 0x30c2 */
            {8'h00}, /* 0x30c1 */
            {8'h00}, /* 0x30c0 */
            {8'h00}, /* 0x30bf */
            {8'h00}, /* 0x30be */
            {8'h00}, /* 0x30bd */
            {8'h00}, /* 0x30bc */
            {8'h00}, /* 0x30bb */
            {8'h00}, /* 0x30ba */
            {8'h00}, /* 0x30b9 */
            {8'h00}, /* 0x30b8 */
            {8'h00}, /* 0x30b7 */
            {8'h00}, /* 0x30b6 */
            {8'h00}, /* 0x30b5 */
            {8'h00}, /* 0x30b4 */
            {8'h00}, /* 0x30b3 */
            {8'h00}, /* 0x30b2 */
            {8'h00}, /* 0x30b1 */
            {8'h00}, /* 0x30b0 */
            {8'h00}, /* 0x30af */
            {8'h00}, /* 0x30ae */
            {8'h00}, /* 0x30ad */
            {8'h00}, /* 0x30ac */
            {8'h00}, /* 0x30ab */
            {8'h00}, /* 0x30aa */
            {8'h00}, /* 0x30a9 */
            {8'h00}, /* 0x30a8 */
            {8'h00}, /* 0x30a7 */
            {8'h00}, /* 0x30a6 */
            {8'h00}, /* 0x30a5 */
            {8'h00}, /* 0x30a4 */
            {8'h00}, /* 0x30a3 */
            {8'h00}, /* 0x30a2 */
            {8'h00}, /* 0x30a1 */
            {8'h00}, /* 0x30a0 */
            {8'h00}, /* 0x309f */
            {8'h00}, /* 0x309e */
            {8'h00}, /* 0x309d */
            {8'h00}, /* 0x309c */
            {8'h00}, /* 0x309b */
            {8'h00}, /* 0x309a */
            {8'h00}, /* 0x3099 */
            {8'h00}, /* 0x3098 */
            {8'h00}, /* 0x3097 */
            {8'h00}, /* 0x3096 */
            {8'h00}, /* 0x3095 */
            {8'h00}, /* 0x3094 */
            {8'h00}, /* 0x3093 */
            {8'h00}, /* 0x3092 */
            {8'h00}, /* 0x3091 */
            {8'h00}, /* 0x3090 */
            {8'h00}, /* 0x308f */
            {8'h00}, /* 0x308e */
            {8'h00}, /* 0x308d */
            {8'h00}, /* 0x308c */
            {8'h00}, /* 0x308b */
            {8'h00}, /* 0x308a */
            {8'h00}, /* 0x3089 */
            {8'h00}, /* 0x3088 */
            {8'h00}, /* 0x3087 */
            {8'h00}, /* 0x3086 */
            {8'h00}, /* 0x3085 */
            {8'h00}, /* 0x3084 */
            {8'h00}, /* 0x3083 */
            {8'h00}, /* 0x3082 */
            {8'h00}, /* 0x3081 */
            {8'h00}, /* 0x3080 */
            {8'h00}, /* 0x307f */
            {8'h00}, /* 0x307e */
            {8'h00}, /* 0x307d */
            {8'h00}, /* 0x307c */
            {8'h00}, /* 0x307b */
            {8'h00}, /* 0x307a */
            {8'h00}, /* 0x3079 */
            {8'h00}, /* 0x3078 */
            {8'h00}, /* 0x3077 */
            {8'h00}, /* 0x3076 */
            {8'h00}, /* 0x3075 */
            {8'h00}, /* 0x3074 */
            {8'h00}, /* 0x3073 */
            {8'h00}, /* 0x3072 */
            {8'h00}, /* 0x3071 */
            {8'h00}, /* 0x3070 */
            {8'h00}, /* 0x306f */
            {8'h00}, /* 0x306e */
            {8'h00}, /* 0x306d */
            {8'h00}, /* 0x306c */
            {8'h00}, /* 0x306b */
            {8'h00}, /* 0x306a */
            {8'h00}, /* 0x3069 */
            {8'h00}, /* 0x3068 */
            {8'h00}, /* 0x3067 */
            {8'h00}, /* 0x3066 */
            {8'h00}, /* 0x3065 */
            {8'h00}, /* 0x3064 */
            {8'h00}, /* 0x3063 */
            {8'h00}, /* 0x3062 */
            {8'h00}, /* 0x3061 */
            {8'h00}, /* 0x3060 */
            {8'h00}, /* 0x305f */
            {8'h00}, /* 0x305e */
            {8'h00}, /* 0x305d */
            {8'h00}, /* 0x305c */
            {8'h00}, /* 0x305b */
            {8'h00}, /* 0x305a */
            {8'h00}, /* 0x3059 */
            {8'h00}, /* 0x3058 */
            {8'h00}, /* 0x3057 */
            {8'h00}, /* 0x3056 */
            {8'h00}, /* 0x3055 */
            {8'h00}, /* 0x3054 */
            {8'h00}, /* 0x3053 */
            {8'h00}, /* 0x3052 */
            {8'h00}, /* 0x3051 */
            {8'h00}, /* 0x3050 */
            {8'h00}, /* 0x304f */
            {8'h00}, /* 0x304e */
            {8'h00}, /* 0x304d */
            {8'h00}, /* 0x304c */
            {8'h00}, /* 0x304b */
            {8'h00}, /* 0x304a */
            {8'h00}, /* 0x3049 */
            {8'h00}, /* 0x3048 */
            {8'h00}, /* 0x3047 */
            {8'h00}, /* 0x3046 */
            {8'h00}, /* 0x3045 */
            {8'h00}, /* 0x3044 */
            {8'h00}, /* 0x3043 */
            {8'h00}, /* 0x3042 */
            {8'h00}, /* 0x3041 */
            {8'h00}, /* 0x3040 */
            {8'h00}, /* 0x303f */
            {8'h00}, /* 0x303e */
            {8'h00}, /* 0x303d */
            {8'h00}, /* 0x303c */
            {8'h00}, /* 0x303b */
            {8'h00}, /* 0x303a */
            {8'h00}, /* 0x3039 */
            {8'h00}, /* 0x3038 */
            {8'h00}, /* 0x3037 */
            {8'h00}, /* 0x3036 */
            {8'h00}, /* 0x3035 */
            {8'h00}, /* 0x3034 */
            {8'h00}, /* 0x3033 */
            {8'h00}, /* 0x3032 */
            {8'h00}, /* 0x3031 */
            {8'h00}, /* 0x3030 */
            {8'h00}, /* 0x302f */
            {8'h00}, /* 0x302e */
            {8'h00}, /* 0x302d */
            {8'h00}, /* 0x302c */
            {8'h00}, /* 0x302b */
            {8'h00}, /* 0x302a */
            {8'h00}, /* 0x3029 */
            {8'h00}, /* 0x3028 */
            {8'h00}, /* 0x3027 */
            {8'h00}, /* 0x3026 */
            {8'h00}, /* 0x3025 */
            {8'h00}, /* 0x3024 */
            {8'h00}, /* 0x3023 */
            {8'h00}, /* 0x3022 */
            {8'h00}, /* 0x3021 */
            {8'h00}, /* 0x3020 */
            {8'h00}, /* 0x301f */
            {8'h00}, /* 0x301e */
            {8'h00}, /* 0x301d */
            {8'h00}, /* 0x301c */
            {8'h00}, /* 0x301b */
            {8'h00}, /* 0x301a */
            {8'h00}, /* 0x3019 */
            {8'h00}, /* 0x3018 */
            {8'h00}, /* 0x3017 */
            {8'h00}, /* 0x3016 */
            {8'h00}, /* 0x3015 */
            {8'h00}, /* 0x3014 */
            {8'h00}, /* 0x3013 */
            {8'h00}, /* 0x3012 */
            {8'h00}, /* 0x3011 */
            {8'h00}, /* 0x3010 */
            {8'h00}, /* 0x300f */
            {8'h00}, /* 0x300e */
            {8'h00}, /* 0x300d */
            {8'h00}, /* 0x300c */
            {8'h00}, /* 0x300b */
            {8'h00}, /* 0x300a */
            {8'h00}, /* 0x3009 */
            {8'h00}, /* 0x3008 */
            {8'h00}, /* 0x3007 */
            {8'h00}, /* 0x3006 */
            {8'h00}, /* 0x3005 */
            {8'h00}, /* 0x3004 */
            {8'h00}, /* 0x3003 */
            {8'h00}, /* 0x3002 */
            {8'h00}, /* 0x3001 */
            {8'h00}, /* 0x3000 */
            {8'h00}, /* 0x2fff */
            {8'h00}, /* 0x2ffe */
            {8'h00}, /* 0x2ffd */
            {8'h00}, /* 0x2ffc */
            {8'h00}, /* 0x2ffb */
            {8'h00}, /* 0x2ffa */
            {8'h00}, /* 0x2ff9 */
            {8'h00}, /* 0x2ff8 */
            {8'h00}, /* 0x2ff7 */
            {8'h00}, /* 0x2ff6 */
            {8'h00}, /* 0x2ff5 */
            {8'h00}, /* 0x2ff4 */
            {8'h00}, /* 0x2ff3 */
            {8'h00}, /* 0x2ff2 */
            {8'h00}, /* 0x2ff1 */
            {8'h00}, /* 0x2ff0 */
            {8'h00}, /* 0x2fef */
            {8'h00}, /* 0x2fee */
            {8'h00}, /* 0x2fed */
            {8'h00}, /* 0x2fec */
            {8'h00}, /* 0x2feb */
            {8'h00}, /* 0x2fea */
            {8'h00}, /* 0x2fe9 */
            {8'h00}, /* 0x2fe8 */
            {8'h00}, /* 0x2fe7 */
            {8'h00}, /* 0x2fe6 */
            {8'h00}, /* 0x2fe5 */
            {8'h00}, /* 0x2fe4 */
            {8'h00}, /* 0x2fe3 */
            {8'h00}, /* 0x2fe2 */
            {8'h00}, /* 0x2fe1 */
            {8'h00}, /* 0x2fe0 */
            {8'h00}, /* 0x2fdf */
            {8'h00}, /* 0x2fde */
            {8'h00}, /* 0x2fdd */
            {8'h00}, /* 0x2fdc */
            {8'h00}, /* 0x2fdb */
            {8'h00}, /* 0x2fda */
            {8'h00}, /* 0x2fd9 */
            {8'h00}, /* 0x2fd8 */
            {8'h00}, /* 0x2fd7 */
            {8'h00}, /* 0x2fd6 */
            {8'h00}, /* 0x2fd5 */
            {8'h00}, /* 0x2fd4 */
            {8'h00}, /* 0x2fd3 */
            {8'h00}, /* 0x2fd2 */
            {8'h00}, /* 0x2fd1 */
            {8'h00}, /* 0x2fd0 */
            {8'h00}, /* 0x2fcf */
            {8'h00}, /* 0x2fce */
            {8'h00}, /* 0x2fcd */
            {8'h00}, /* 0x2fcc */
            {8'h00}, /* 0x2fcb */
            {8'h00}, /* 0x2fca */
            {8'h00}, /* 0x2fc9 */
            {8'h00}, /* 0x2fc8 */
            {8'h00}, /* 0x2fc7 */
            {8'h00}, /* 0x2fc6 */
            {8'h00}, /* 0x2fc5 */
            {8'h00}, /* 0x2fc4 */
            {8'h00}, /* 0x2fc3 */
            {8'h00}, /* 0x2fc2 */
            {8'h00}, /* 0x2fc1 */
            {8'h00}, /* 0x2fc0 */
            {8'h00}, /* 0x2fbf */
            {8'h00}, /* 0x2fbe */
            {8'h00}, /* 0x2fbd */
            {8'h00}, /* 0x2fbc */
            {8'h00}, /* 0x2fbb */
            {8'h00}, /* 0x2fba */
            {8'h00}, /* 0x2fb9 */
            {8'h00}, /* 0x2fb8 */
            {8'h00}, /* 0x2fb7 */
            {8'h00}, /* 0x2fb6 */
            {8'h00}, /* 0x2fb5 */
            {8'h00}, /* 0x2fb4 */
            {8'h00}, /* 0x2fb3 */
            {8'h00}, /* 0x2fb2 */
            {8'h00}, /* 0x2fb1 */
            {8'h00}, /* 0x2fb0 */
            {8'h00}, /* 0x2faf */
            {8'h00}, /* 0x2fae */
            {8'h00}, /* 0x2fad */
            {8'h00}, /* 0x2fac */
            {8'h00}, /* 0x2fab */
            {8'h00}, /* 0x2faa */
            {8'h00}, /* 0x2fa9 */
            {8'h00}, /* 0x2fa8 */
            {8'h00}, /* 0x2fa7 */
            {8'h00}, /* 0x2fa6 */
            {8'h00}, /* 0x2fa5 */
            {8'h00}, /* 0x2fa4 */
            {8'h00}, /* 0x2fa3 */
            {8'h00}, /* 0x2fa2 */
            {8'h00}, /* 0x2fa1 */
            {8'h00}, /* 0x2fa0 */
            {8'h00}, /* 0x2f9f */
            {8'h00}, /* 0x2f9e */
            {8'h00}, /* 0x2f9d */
            {8'h00}, /* 0x2f9c */
            {8'h00}, /* 0x2f9b */
            {8'h00}, /* 0x2f9a */
            {8'h00}, /* 0x2f99 */
            {8'h00}, /* 0x2f98 */
            {8'h00}, /* 0x2f97 */
            {8'h00}, /* 0x2f96 */
            {8'h00}, /* 0x2f95 */
            {8'h00}, /* 0x2f94 */
            {8'h00}, /* 0x2f93 */
            {8'h00}, /* 0x2f92 */
            {8'h00}, /* 0x2f91 */
            {8'h00}, /* 0x2f90 */
            {8'h00}, /* 0x2f8f */
            {8'h00}, /* 0x2f8e */
            {8'h00}, /* 0x2f8d */
            {8'h00}, /* 0x2f8c */
            {8'h00}, /* 0x2f8b */
            {8'h00}, /* 0x2f8a */
            {8'h00}, /* 0x2f89 */
            {8'h00}, /* 0x2f88 */
            {8'h00}, /* 0x2f87 */
            {8'h00}, /* 0x2f86 */
            {8'h00}, /* 0x2f85 */
            {8'h00}, /* 0x2f84 */
            {8'h00}, /* 0x2f83 */
            {8'h00}, /* 0x2f82 */
            {8'h00}, /* 0x2f81 */
            {8'h00}, /* 0x2f80 */
            {8'h00}, /* 0x2f7f */
            {8'h00}, /* 0x2f7e */
            {8'h00}, /* 0x2f7d */
            {8'h00}, /* 0x2f7c */
            {8'h00}, /* 0x2f7b */
            {8'h00}, /* 0x2f7a */
            {8'h00}, /* 0x2f79 */
            {8'h00}, /* 0x2f78 */
            {8'h00}, /* 0x2f77 */
            {8'h00}, /* 0x2f76 */
            {8'h00}, /* 0x2f75 */
            {8'h00}, /* 0x2f74 */
            {8'h00}, /* 0x2f73 */
            {8'h00}, /* 0x2f72 */
            {8'h00}, /* 0x2f71 */
            {8'h00}, /* 0x2f70 */
            {8'h00}, /* 0x2f6f */
            {8'h00}, /* 0x2f6e */
            {8'h00}, /* 0x2f6d */
            {8'h00}, /* 0x2f6c */
            {8'h00}, /* 0x2f6b */
            {8'h00}, /* 0x2f6a */
            {8'h00}, /* 0x2f69 */
            {8'h00}, /* 0x2f68 */
            {8'h00}, /* 0x2f67 */
            {8'h00}, /* 0x2f66 */
            {8'h00}, /* 0x2f65 */
            {8'h00}, /* 0x2f64 */
            {8'h00}, /* 0x2f63 */
            {8'h00}, /* 0x2f62 */
            {8'h00}, /* 0x2f61 */
            {8'h00}, /* 0x2f60 */
            {8'h00}, /* 0x2f5f */
            {8'h00}, /* 0x2f5e */
            {8'h00}, /* 0x2f5d */
            {8'h00}, /* 0x2f5c */
            {8'h00}, /* 0x2f5b */
            {8'h00}, /* 0x2f5a */
            {8'h00}, /* 0x2f59 */
            {8'h00}, /* 0x2f58 */
            {8'h00}, /* 0x2f57 */
            {8'h00}, /* 0x2f56 */
            {8'h00}, /* 0x2f55 */
            {8'h00}, /* 0x2f54 */
            {8'h00}, /* 0x2f53 */
            {8'h00}, /* 0x2f52 */
            {8'h00}, /* 0x2f51 */
            {8'h00}, /* 0x2f50 */
            {8'h00}, /* 0x2f4f */
            {8'h00}, /* 0x2f4e */
            {8'h00}, /* 0x2f4d */
            {8'h00}, /* 0x2f4c */
            {8'h00}, /* 0x2f4b */
            {8'h00}, /* 0x2f4a */
            {8'h00}, /* 0x2f49 */
            {8'h00}, /* 0x2f48 */
            {8'h00}, /* 0x2f47 */
            {8'h00}, /* 0x2f46 */
            {8'h00}, /* 0x2f45 */
            {8'h00}, /* 0x2f44 */
            {8'h00}, /* 0x2f43 */
            {8'h00}, /* 0x2f42 */
            {8'h00}, /* 0x2f41 */
            {8'h00}, /* 0x2f40 */
            {8'h00}, /* 0x2f3f */
            {8'h00}, /* 0x2f3e */
            {8'h00}, /* 0x2f3d */
            {8'h00}, /* 0x2f3c */
            {8'h00}, /* 0x2f3b */
            {8'h00}, /* 0x2f3a */
            {8'h00}, /* 0x2f39 */
            {8'h00}, /* 0x2f38 */
            {8'h00}, /* 0x2f37 */
            {8'h00}, /* 0x2f36 */
            {8'h00}, /* 0x2f35 */
            {8'h00}, /* 0x2f34 */
            {8'h00}, /* 0x2f33 */
            {8'h00}, /* 0x2f32 */
            {8'h00}, /* 0x2f31 */
            {8'h00}, /* 0x2f30 */
            {8'h00}, /* 0x2f2f */
            {8'h00}, /* 0x2f2e */
            {8'h00}, /* 0x2f2d */
            {8'h00}, /* 0x2f2c */
            {8'h00}, /* 0x2f2b */
            {8'h00}, /* 0x2f2a */
            {8'h00}, /* 0x2f29 */
            {8'h00}, /* 0x2f28 */
            {8'h00}, /* 0x2f27 */
            {8'h00}, /* 0x2f26 */
            {8'h00}, /* 0x2f25 */
            {8'h00}, /* 0x2f24 */
            {8'h00}, /* 0x2f23 */
            {8'h00}, /* 0x2f22 */
            {8'h00}, /* 0x2f21 */
            {8'h00}, /* 0x2f20 */
            {8'h00}, /* 0x2f1f */
            {8'h00}, /* 0x2f1e */
            {8'h00}, /* 0x2f1d */
            {8'h00}, /* 0x2f1c */
            {8'h00}, /* 0x2f1b */
            {8'h00}, /* 0x2f1a */
            {8'h00}, /* 0x2f19 */
            {8'h00}, /* 0x2f18 */
            {8'h00}, /* 0x2f17 */
            {8'h00}, /* 0x2f16 */
            {8'h00}, /* 0x2f15 */
            {8'h00}, /* 0x2f14 */
            {8'h00}, /* 0x2f13 */
            {8'h00}, /* 0x2f12 */
            {8'h00}, /* 0x2f11 */
            {8'h00}, /* 0x2f10 */
            {8'h00}, /* 0x2f0f */
            {8'h00}, /* 0x2f0e */
            {8'h00}, /* 0x2f0d */
            {8'h00}, /* 0x2f0c */
            {8'h00}, /* 0x2f0b */
            {8'h00}, /* 0x2f0a */
            {8'h00}, /* 0x2f09 */
            {8'h00}, /* 0x2f08 */
            {8'h00}, /* 0x2f07 */
            {8'h00}, /* 0x2f06 */
            {8'h00}, /* 0x2f05 */
            {8'h00}, /* 0x2f04 */
            {8'h00}, /* 0x2f03 */
            {8'h00}, /* 0x2f02 */
            {8'h00}, /* 0x2f01 */
            {8'h00}, /* 0x2f00 */
            {8'h00}, /* 0x2eff */
            {8'h00}, /* 0x2efe */
            {8'h00}, /* 0x2efd */
            {8'h00}, /* 0x2efc */
            {8'h00}, /* 0x2efb */
            {8'h00}, /* 0x2efa */
            {8'h00}, /* 0x2ef9 */
            {8'h00}, /* 0x2ef8 */
            {8'h00}, /* 0x2ef7 */
            {8'h00}, /* 0x2ef6 */
            {8'h00}, /* 0x2ef5 */
            {8'h00}, /* 0x2ef4 */
            {8'h00}, /* 0x2ef3 */
            {8'h00}, /* 0x2ef2 */
            {8'h00}, /* 0x2ef1 */
            {8'h00}, /* 0x2ef0 */
            {8'h00}, /* 0x2eef */
            {8'h00}, /* 0x2eee */
            {8'h00}, /* 0x2eed */
            {8'h00}, /* 0x2eec */
            {8'h00}, /* 0x2eeb */
            {8'h00}, /* 0x2eea */
            {8'h00}, /* 0x2ee9 */
            {8'h00}, /* 0x2ee8 */
            {8'h00}, /* 0x2ee7 */
            {8'h00}, /* 0x2ee6 */
            {8'h00}, /* 0x2ee5 */
            {8'h00}, /* 0x2ee4 */
            {8'h00}, /* 0x2ee3 */
            {8'h00}, /* 0x2ee2 */
            {8'h00}, /* 0x2ee1 */
            {8'h00}, /* 0x2ee0 */
            {8'h00}, /* 0x2edf */
            {8'h00}, /* 0x2ede */
            {8'h00}, /* 0x2edd */
            {8'h00}, /* 0x2edc */
            {8'h00}, /* 0x2edb */
            {8'h00}, /* 0x2eda */
            {8'h00}, /* 0x2ed9 */
            {8'h00}, /* 0x2ed8 */
            {8'h00}, /* 0x2ed7 */
            {8'h00}, /* 0x2ed6 */
            {8'h00}, /* 0x2ed5 */
            {8'h00}, /* 0x2ed4 */
            {8'h00}, /* 0x2ed3 */
            {8'h00}, /* 0x2ed2 */
            {8'h00}, /* 0x2ed1 */
            {8'h00}, /* 0x2ed0 */
            {8'h00}, /* 0x2ecf */
            {8'h00}, /* 0x2ece */
            {8'h00}, /* 0x2ecd */
            {8'h00}, /* 0x2ecc */
            {8'h00}, /* 0x2ecb */
            {8'h00}, /* 0x2eca */
            {8'h00}, /* 0x2ec9 */
            {8'h00}, /* 0x2ec8 */
            {8'h00}, /* 0x2ec7 */
            {8'h00}, /* 0x2ec6 */
            {8'h00}, /* 0x2ec5 */
            {8'h00}, /* 0x2ec4 */
            {8'h00}, /* 0x2ec3 */
            {8'h00}, /* 0x2ec2 */
            {8'h00}, /* 0x2ec1 */
            {8'h00}, /* 0x2ec0 */
            {8'h00}, /* 0x2ebf */
            {8'h00}, /* 0x2ebe */
            {8'h00}, /* 0x2ebd */
            {8'h00}, /* 0x2ebc */
            {8'h00}, /* 0x2ebb */
            {8'h00}, /* 0x2eba */
            {8'h00}, /* 0x2eb9 */
            {8'h00}, /* 0x2eb8 */
            {8'h00}, /* 0x2eb7 */
            {8'h00}, /* 0x2eb6 */
            {8'h00}, /* 0x2eb5 */
            {8'h00}, /* 0x2eb4 */
            {8'h00}, /* 0x2eb3 */
            {8'h00}, /* 0x2eb2 */
            {8'h00}, /* 0x2eb1 */
            {8'h00}, /* 0x2eb0 */
            {8'h00}, /* 0x2eaf */
            {8'h00}, /* 0x2eae */
            {8'h00}, /* 0x2ead */
            {8'h00}, /* 0x2eac */
            {8'h00}, /* 0x2eab */
            {8'h00}, /* 0x2eaa */
            {8'h00}, /* 0x2ea9 */
            {8'h00}, /* 0x2ea8 */
            {8'h00}, /* 0x2ea7 */
            {8'h00}, /* 0x2ea6 */
            {8'h00}, /* 0x2ea5 */
            {8'h00}, /* 0x2ea4 */
            {8'h00}, /* 0x2ea3 */
            {8'h00}, /* 0x2ea2 */
            {8'h00}, /* 0x2ea1 */
            {8'h00}, /* 0x2ea0 */
            {8'h00}, /* 0x2e9f */
            {8'h00}, /* 0x2e9e */
            {8'h00}, /* 0x2e9d */
            {8'h00}, /* 0x2e9c */
            {8'h00}, /* 0x2e9b */
            {8'h00}, /* 0x2e9a */
            {8'h00}, /* 0x2e99 */
            {8'h00}, /* 0x2e98 */
            {8'h00}, /* 0x2e97 */
            {8'h00}, /* 0x2e96 */
            {8'h00}, /* 0x2e95 */
            {8'h00}, /* 0x2e94 */
            {8'h00}, /* 0x2e93 */
            {8'h00}, /* 0x2e92 */
            {8'h00}, /* 0x2e91 */
            {8'h00}, /* 0x2e90 */
            {8'h00}, /* 0x2e8f */
            {8'h00}, /* 0x2e8e */
            {8'h00}, /* 0x2e8d */
            {8'h00}, /* 0x2e8c */
            {8'h00}, /* 0x2e8b */
            {8'h00}, /* 0x2e8a */
            {8'h00}, /* 0x2e89 */
            {8'h00}, /* 0x2e88 */
            {8'h00}, /* 0x2e87 */
            {8'h00}, /* 0x2e86 */
            {8'h00}, /* 0x2e85 */
            {8'h00}, /* 0x2e84 */
            {8'h00}, /* 0x2e83 */
            {8'h00}, /* 0x2e82 */
            {8'h00}, /* 0x2e81 */
            {8'h00}, /* 0x2e80 */
            {8'h00}, /* 0x2e7f */
            {8'h00}, /* 0x2e7e */
            {8'h00}, /* 0x2e7d */
            {8'h00}, /* 0x2e7c */
            {8'h00}, /* 0x2e7b */
            {8'h00}, /* 0x2e7a */
            {8'h00}, /* 0x2e79 */
            {8'h00}, /* 0x2e78 */
            {8'h00}, /* 0x2e77 */
            {8'h00}, /* 0x2e76 */
            {8'h00}, /* 0x2e75 */
            {8'h00}, /* 0x2e74 */
            {8'h00}, /* 0x2e73 */
            {8'h00}, /* 0x2e72 */
            {8'h00}, /* 0x2e71 */
            {8'h00}, /* 0x2e70 */
            {8'h00}, /* 0x2e6f */
            {8'h00}, /* 0x2e6e */
            {8'h00}, /* 0x2e6d */
            {8'h00}, /* 0x2e6c */
            {8'h00}, /* 0x2e6b */
            {8'h00}, /* 0x2e6a */
            {8'h00}, /* 0x2e69 */
            {8'h00}, /* 0x2e68 */
            {8'h00}, /* 0x2e67 */
            {8'h00}, /* 0x2e66 */
            {8'h00}, /* 0x2e65 */
            {8'h00}, /* 0x2e64 */
            {8'h00}, /* 0x2e63 */
            {8'h00}, /* 0x2e62 */
            {8'h00}, /* 0x2e61 */
            {8'h00}, /* 0x2e60 */
            {8'h00}, /* 0x2e5f */
            {8'h00}, /* 0x2e5e */
            {8'h00}, /* 0x2e5d */
            {8'h00}, /* 0x2e5c */
            {8'h00}, /* 0x2e5b */
            {8'h00}, /* 0x2e5a */
            {8'h00}, /* 0x2e59 */
            {8'h00}, /* 0x2e58 */
            {8'h00}, /* 0x2e57 */
            {8'h00}, /* 0x2e56 */
            {8'h00}, /* 0x2e55 */
            {8'h00}, /* 0x2e54 */
            {8'h00}, /* 0x2e53 */
            {8'h00}, /* 0x2e52 */
            {8'h00}, /* 0x2e51 */
            {8'h00}, /* 0x2e50 */
            {8'h00}, /* 0x2e4f */
            {8'h00}, /* 0x2e4e */
            {8'h00}, /* 0x2e4d */
            {8'h00}, /* 0x2e4c */
            {8'h00}, /* 0x2e4b */
            {8'h00}, /* 0x2e4a */
            {8'h00}, /* 0x2e49 */
            {8'h00}, /* 0x2e48 */
            {8'h00}, /* 0x2e47 */
            {8'h00}, /* 0x2e46 */
            {8'h00}, /* 0x2e45 */
            {8'h00}, /* 0x2e44 */
            {8'h00}, /* 0x2e43 */
            {8'h00}, /* 0x2e42 */
            {8'h00}, /* 0x2e41 */
            {8'h00}, /* 0x2e40 */
            {8'h00}, /* 0x2e3f */
            {8'h00}, /* 0x2e3e */
            {8'h00}, /* 0x2e3d */
            {8'h00}, /* 0x2e3c */
            {8'h00}, /* 0x2e3b */
            {8'h00}, /* 0x2e3a */
            {8'h00}, /* 0x2e39 */
            {8'h00}, /* 0x2e38 */
            {8'h00}, /* 0x2e37 */
            {8'h00}, /* 0x2e36 */
            {8'h00}, /* 0x2e35 */
            {8'h00}, /* 0x2e34 */
            {8'h00}, /* 0x2e33 */
            {8'h00}, /* 0x2e32 */
            {8'h00}, /* 0x2e31 */
            {8'h00}, /* 0x2e30 */
            {8'h00}, /* 0x2e2f */
            {8'h00}, /* 0x2e2e */
            {8'h00}, /* 0x2e2d */
            {8'h00}, /* 0x2e2c */
            {8'h00}, /* 0x2e2b */
            {8'h00}, /* 0x2e2a */
            {8'h00}, /* 0x2e29 */
            {8'h00}, /* 0x2e28 */
            {8'h00}, /* 0x2e27 */
            {8'h00}, /* 0x2e26 */
            {8'h00}, /* 0x2e25 */
            {8'h00}, /* 0x2e24 */
            {8'h00}, /* 0x2e23 */
            {8'h00}, /* 0x2e22 */
            {8'h00}, /* 0x2e21 */
            {8'h00}, /* 0x2e20 */
            {8'h00}, /* 0x2e1f */
            {8'h00}, /* 0x2e1e */
            {8'h00}, /* 0x2e1d */
            {8'h00}, /* 0x2e1c */
            {8'h00}, /* 0x2e1b */
            {8'h00}, /* 0x2e1a */
            {8'h00}, /* 0x2e19 */
            {8'h00}, /* 0x2e18 */
            {8'h00}, /* 0x2e17 */
            {8'h00}, /* 0x2e16 */
            {8'h00}, /* 0x2e15 */
            {8'h00}, /* 0x2e14 */
            {8'h00}, /* 0x2e13 */
            {8'h00}, /* 0x2e12 */
            {8'h00}, /* 0x2e11 */
            {8'h00}, /* 0x2e10 */
            {8'h00}, /* 0x2e0f */
            {8'h00}, /* 0x2e0e */
            {8'h00}, /* 0x2e0d */
            {8'h00}, /* 0x2e0c */
            {8'h00}, /* 0x2e0b */
            {8'h00}, /* 0x2e0a */
            {8'h00}, /* 0x2e09 */
            {8'h00}, /* 0x2e08 */
            {8'h00}, /* 0x2e07 */
            {8'h00}, /* 0x2e06 */
            {8'h00}, /* 0x2e05 */
            {8'h00}, /* 0x2e04 */
            {8'h00}, /* 0x2e03 */
            {8'h00}, /* 0x2e02 */
            {8'h00}, /* 0x2e01 */
            {8'h00}, /* 0x2e00 */
            {8'h00}, /* 0x2dff */
            {8'h00}, /* 0x2dfe */
            {8'h00}, /* 0x2dfd */
            {8'h00}, /* 0x2dfc */
            {8'h00}, /* 0x2dfb */
            {8'h00}, /* 0x2dfa */
            {8'h00}, /* 0x2df9 */
            {8'h00}, /* 0x2df8 */
            {8'h00}, /* 0x2df7 */
            {8'h00}, /* 0x2df6 */
            {8'h00}, /* 0x2df5 */
            {8'h00}, /* 0x2df4 */
            {8'h00}, /* 0x2df3 */
            {8'h00}, /* 0x2df2 */
            {8'h00}, /* 0x2df1 */
            {8'h00}, /* 0x2df0 */
            {8'h00}, /* 0x2def */
            {8'h00}, /* 0x2dee */
            {8'h00}, /* 0x2ded */
            {8'h00}, /* 0x2dec */
            {8'h00}, /* 0x2deb */
            {8'h00}, /* 0x2dea */
            {8'h00}, /* 0x2de9 */
            {8'h00}, /* 0x2de8 */
            {8'h00}, /* 0x2de7 */
            {8'h00}, /* 0x2de6 */
            {8'h00}, /* 0x2de5 */
            {8'h00}, /* 0x2de4 */
            {8'h00}, /* 0x2de3 */
            {8'h00}, /* 0x2de2 */
            {8'h00}, /* 0x2de1 */
            {8'h00}, /* 0x2de0 */
            {8'h00}, /* 0x2ddf */
            {8'h00}, /* 0x2dde */
            {8'h00}, /* 0x2ddd */
            {8'h00}, /* 0x2ddc */
            {8'h00}, /* 0x2ddb */
            {8'h00}, /* 0x2dda */
            {8'h00}, /* 0x2dd9 */
            {8'h00}, /* 0x2dd8 */
            {8'h00}, /* 0x2dd7 */
            {8'h00}, /* 0x2dd6 */
            {8'h00}, /* 0x2dd5 */
            {8'h00}, /* 0x2dd4 */
            {8'h00}, /* 0x2dd3 */
            {8'h00}, /* 0x2dd2 */
            {8'h00}, /* 0x2dd1 */
            {8'h00}, /* 0x2dd0 */
            {8'h00}, /* 0x2dcf */
            {8'h00}, /* 0x2dce */
            {8'h00}, /* 0x2dcd */
            {8'h00}, /* 0x2dcc */
            {8'h00}, /* 0x2dcb */
            {8'h00}, /* 0x2dca */
            {8'h00}, /* 0x2dc9 */
            {8'h00}, /* 0x2dc8 */
            {8'h00}, /* 0x2dc7 */
            {8'h00}, /* 0x2dc6 */
            {8'h00}, /* 0x2dc5 */
            {8'h00}, /* 0x2dc4 */
            {8'h00}, /* 0x2dc3 */
            {8'h00}, /* 0x2dc2 */
            {8'h00}, /* 0x2dc1 */
            {8'h00}, /* 0x2dc0 */
            {8'h00}, /* 0x2dbf */
            {8'h00}, /* 0x2dbe */
            {8'h00}, /* 0x2dbd */
            {8'h00}, /* 0x2dbc */
            {8'h00}, /* 0x2dbb */
            {8'h00}, /* 0x2dba */
            {8'h00}, /* 0x2db9 */
            {8'h00}, /* 0x2db8 */
            {8'h00}, /* 0x2db7 */
            {8'h00}, /* 0x2db6 */
            {8'h00}, /* 0x2db5 */
            {8'h00}, /* 0x2db4 */
            {8'h00}, /* 0x2db3 */
            {8'h00}, /* 0x2db2 */
            {8'h00}, /* 0x2db1 */
            {8'h00}, /* 0x2db0 */
            {8'h00}, /* 0x2daf */
            {8'h00}, /* 0x2dae */
            {8'h00}, /* 0x2dad */
            {8'h00}, /* 0x2dac */
            {8'h00}, /* 0x2dab */
            {8'h00}, /* 0x2daa */
            {8'h00}, /* 0x2da9 */
            {8'h00}, /* 0x2da8 */
            {8'h00}, /* 0x2da7 */
            {8'h00}, /* 0x2da6 */
            {8'h00}, /* 0x2da5 */
            {8'h00}, /* 0x2da4 */
            {8'h00}, /* 0x2da3 */
            {8'h00}, /* 0x2da2 */
            {8'h00}, /* 0x2da1 */
            {8'h00}, /* 0x2da0 */
            {8'h00}, /* 0x2d9f */
            {8'h00}, /* 0x2d9e */
            {8'h00}, /* 0x2d9d */
            {8'h00}, /* 0x2d9c */
            {8'h00}, /* 0x2d9b */
            {8'h00}, /* 0x2d9a */
            {8'h00}, /* 0x2d99 */
            {8'h00}, /* 0x2d98 */
            {8'h00}, /* 0x2d97 */
            {8'h00}, /* 0x2d96 */
            {8'h00}, /* 0x2d95 */
            {8'h00}, /* 0x2d94 */
            {8'h00}, /* 0x2d93 */
            {8'h00}, /* 0x2d92 */
            {8'h00}, /* 0x2d91 */
            {8'h00}, /* 0x2d90 */
            {8'h00}, /* 0x2d8f */
            {8'h00}, /* 0x2d8e */
            {8'h00}, /* 0x2d8d */
            {8'h00}, /* 0x2d8c */
            {8'h00}, /* 0x2d8b */
            {8'h00}, /* 0x2d8a */
            {8'h00}, /* 0x2d89 */
            {8'h00}, /* 0x2d88 */
            {8'h00}, /* 0x2d87 */
            {8'h00}, /* 0x2d86 */
            {8'h00}, /* 0x2d85 */
            {8'h00}, /* 0x2d84 */
            {8'h00}, /* 0x2d83 */
            {8'h00}, /* 0x2d82 */
            {8'h00}, /* 0x2d81 */
            {8'h00}, /* 0x2d80 */
            {8'h00}, /* 0x2d7f */
            {8'h00}, /* 0x2d7e */
            {8'h00}, /* 0x2d7d */
            {8'h00}, /* 0x2d7c */
            {8'h00}, /* 0x2d7b */
            {8'h00}, /* 0x2d7a */
            {8'h00}, /* 0x2d79 */
            {8'h00}, /* 0x2d78 */
            {8'h00}, /* 0x2d77 */
            {8'h00}, /* 0x2d76 */
            {8'h00}, /* 0x2d75 */
            {8'h00}, /* 0x2d74 */
            {8'h00}, /* 0x2d73 */
            {8'h00}, /* 0x2d72 */
            {8'h00}, /* 0x2d71 */
            {8'h00}, /* 0x2d70 */
            {8'h00}, /* 0x2d6f */
            {8'h00}, /* 0x2d6e */
            {8'h00}, /* 0x2d6d */
            {8'h00}, /* 0x2d6c */
            {8'h00}, /* 0x2d6b */
            {8'h00}, /* 0x2d6a */
            {8'h00}, /* 0x2d69 */
            {8'h00}, /* 0x2d68 */
            {8'h00}, /* 0x2d67 */
            {8'h00}, /* 0x2d66 */
            {8'h00}, /* 0x2d65 */
            {8'h00}, /* 0x2d64 */
            {8'h00}, /* 0x2d63 */
            {8'h00}, /* 0x2d62 */
            {8'h00}, /* 0x2d61 */
            {8'h00}, /* 0x2d60 */
            {8'h00}, /* 0x2d5f */
            {8'h00}, /* 0x2d5e */
            {8'h00}, /* 0x2d5d */
            {8'h00}, /* 0x2d5c */
            {8'h00}, /* 0x2d5b */
            {8'h00}, /* 0x2d5a */
            {8'h00}, /* 0x2d59 */
            {8'h00}, /* 0x2d58 */
            {8'h00}, /* 0x2d57 */
            {8'h00}, /* 0x2d56 */
            {8'h00}, /* 0x2d55 */
            {8'h00}, /* 0x2d54 */
            {8'h00}, /* 0x2d53 */
            {8'h00}, /* 0x2d52 */
            {8'h00}, /* 0x2d51 */
            {8'h00}, /* 0x2d50 */
            {8'h00}, /* 0x2d4f */
            {8'h00}, /* 0x2d4e */
            {8'h00}, /* 0x2d4d */
            {8'h00}, /* 0x2d4c */
            {8'h00}, /* 0x2d4b */
            {8'h00}, /* 0x2d4a */
            {8'h00}, /* 0x2d49 */
            {8'h00}, /* 0x2d48 */
            {8'h00}, /* 0x2d47 */
            {8'h00}, /* 0x2d46 */
            {8'h00}, /* 0x2d45 */
            {8'h00}, /* 0x2d44 */
            {8'h00}, /* 0x2d43 */
            {8'h00}, /* 0x2d42 */
            {8'h00}, /* 0x2d41 */
            {8'h00}, /* 0x2d40 */
            {8'h00}, /* 0x2d3f */
            {8'h00}, /* 0x2d3e */
            {8'h00}, /* 0x2d3d */
            {8'h00}, /* 0x2d3c */
            {8'h00}, /* 0x2d3b */
            {8'h00}, /* 0x2d3a */
            {8'h00}, /* 0x2d39 */
            {8'h00}, /* 0x2d38 */
            {8'h00}, /* 0x2d37 */
            {8'h00}, /* 0x2d36 */
            {8'h00}, /* 0x2d35 */
            {8'h00}, /* 0x2d34 */
            {8'h00}, /* 0x2d33 */
            {8'h00}, /* 0x2d32 */
            {8'h00}, /* 0x2d31 */
            {8'h00}, /* 0x2d30 */
            {8'h00}, /* 0x2d2f */
            {8'h00}, /* 0x2d2e */
            {8'h00}, /* 0x2d2d */
            {8'h00}, /* 0x2d2c */
            {8'h00}, /* 0x2d2b */
            {8'h00}, /* 0x2d2a */
            {8'h00}, /* 0x2d29 */
            {8'h00}, /* 0x2d28 */
            {8'h00}, /* 0x2d27 */
            {8'h00}, /* 0x2d26 */
            {8'h00}, /* 0x2d25 */
            {8'h00}, /* 0x2d24 */
            {8'h00}, /* 0x2d23 */
            {8'h00}, /* 0x2d22 */
            {8'h00}, /* 0x2d21 */
            {8'h00}, /* 0x2d20 */
            {8'h00}, /* 0x2d1f */
            {8'h00}, /* 0x2d1e */
            {8'h00}, /* 0x2d1d */
            {8'h00}, /* 0x2d1c */
            {8'h00}, /* 0x2d1b */
            {8'h00}, /* 0x2d1a */
            {8'h00}, /* 0x2d19 */
            {8'h00}, /* 0x2d18 */
            {8'h00}, /* 0x2d17 */
            {8'h00}, /* 0x2d16 */
            {8'h00}, /* 0x2d15 */
            {8'h00}, /* 0x2d14 */
            {8'h00}, /* 0x2d13 */
            {8'h00}, /* 0x2d12 */
            {8'h00}, /* 0x2d11 */
            {8'h00}, /* 0x2d10 */
            {8'h00}, /* 0x2d0f */
            {8'h00}, /* 0x2d0e */
            {8'h00}, /* 0x2d0d */
            {8'h00}, /* 0x2d0c */
            {8'h00}, /* 0x2d0b */
            {8'h00}, /* 0x2d0a */
            {8'h00}, /* 0x2d09 */
            {8'h00}, /* 0x2d08 */
            {8'h00}, /* 0x2d07 */
            {8'h00}, /* 0x2d06 */
            {8'h00}, /* 0x2d05 */
            {8'h00}, /* 0x2d04 */
            {8'h00}, /* 0x2d03 */
            {8'h00}, /* 0x2d02 */
            {8'h00}, /* 0x2d01 */
            {8'h00}, /* 0x2d00 */
            {8'h00}, /* 0x2cff */
            {8'h00}, /* 0x2cfe */
            {8'h00}, /* 0x2cfd */
            {8'h00}, /* 0x2cfc */
            {8'h00}, /* 0x2cfb */
            {8'h00}, /* 0x2cfa */
            {8'h00}, /* 0x2cf9 */
            {8'h00}, /* 0x2cf8 */
            {8'h00}, /* 0x2cf7 */
            {8'h00}, /* 0x2cf6 */
            {8'h00}, /* 0x2cf5 */
            {8'h00}, /* 0x2cf4 */
            {8'h00}, /* 0x2cf3 */
            {8'h00}, /* 0x2cf2 */
            {8'h00}, /* 0x2cf1 */
            {8'h00}, /* 0x2cf0 */
            {8'h00}, /* 0x2cef */
            {8'h00}, /* 0x2cee */
            {8'h00}, /* 0x2ced */
            {8'h00}, /* 0x2cec */
            {8'h00}, /* 0x2ceb */
            {8'h00}, /* 0x2cea */
            {8'h00}, /* 0x2ce9 */
            {8'h00}, /* 0x2ce8 */
            {8'h00}, /* 0x2ce7 */
            {8'h00}, /* 0x2ce6 */
            {8'h00}, /* 0x2ce5 */
            {8'h00}, /* 0x2ce4 */
            {8'h00}, /* 0x2ce3 */
            {8'h00}, /* 0x2ce2 */
            {8'h00}, /* 0x2ce1 */
            {8'h00}, /* 0x2ce0 */
            {8'h00}, /* 0x2cdf */
            {8'h00}, /* 0x2cde */
            {8'h00}, /* 0x2cdd */
            {8'h00}, /* 0x2cdc */
            {8'h00}, /* 0x2cdb */
            {8'h00}, /* 0x2cda */
            {8'h00}, /* 0x2cd9 */
            {8'h00}, /* 0x2cd8 */
            {8'h00}, /* 0x2cd7 */
            {8'h00}, /* 0x2cd6 */
            {8'h00}, /* 0x2cd5 */
            {8'h00}, /* 0x2cd4 */
            {8'h00}, /* 0x2cd3 */
            {8'h00}, /* 0x2cd2 */
            {8'h00}, /* 0x2cd1 */
            {8'h00}, /* 0x2cd0 */
            {8'h00}, /* 0x2ccf */
            {8'h00}, /* 0x2cce */
            {8'h00}, /* 0x2ccd */
            {8'h00}, /* 0x2ccc */
            {8'h00}, /* 0x2ccb */
            {8'h00}, /* 0x2cca */
            {8'h00}, /* 0x2cc9 */
            {8'h00}, /* 0x2cc8 */
            {8'h00}, /* 0x2cc7 */
            {8'h00}, /* 0x2cc6 */
            {8'h00}, /* 0x2cc5 */
            {8'h00}, /* 0x2cc4 */
            {8'h00}, /* 0x2cc3 */
            {8'h00}, /* 0x2cc2 */
            {8'h00}, /* 0x2cc1 */
            {8'h00}, /* 0x2cc0 */
            {8'h00}, /* 0x2cbf */
            {8'h00}, /* 0x2cbe */
            {8'h00}, /* 0x2cbd */
            {8'h00}, /* 0x2cbc */
            {8'h00}, /* 0x2cbb */
            {8'h00}, /* 0x2cba */
            {8'h00}, /* 0x2cb9 */
            {8'h00}, /* 0x2cb8 */
            {8'h00}, /* 0x2cb7 */
            {8'h00}, /* 0x2cb6 */
            {8'h00}, /* 0x2cb5 */
            {8'h00}, /* 0x2cb4 */
            {8'h00}, /* 0x2cb3 */
            {8'h00}, /* 0x2cb2 */
            {8'h00}, /* 0x2cb1 */
            {8'h00}, /* 0x2cb0 */
            {8'h00}, /* 0x2caf */
            {8'h00}, /* 0x2cae */
            {8'h00}, /* 0x2cad */
            {8'h00}, /* 0x2cac */
            {8'h00}, /* 0x2cab */
            {8'h00}, /* 0x2caa */
            {8'h00}, /* 0x2ca9 */
            {8'h00}, /* 0x2ca8 */
            {8'h00}, /* 0x2ca7 */
            {8'h00}, /* 0x2ca6 */
            {8'h00}, /* 0x2ca5 */
            {8'h00}, /* 0x2ca4 */
            {8'h00}, /* 0x2ca3 */
            {8'h00}, /* 0x2ca2 */
            {8'h00}, /* 0x2ca1 */
            {8'h00}, /* 0x2ca0 */
            {8'h00}, /* 0x2c9f */
            {8'h00}, /* 0x2c9e */
            {8'h00}, /* 0x2c9d */
            {8'h00}, /* 0x2c9c */
            {8'h00}, /* 0x2c9b */
            {8'h00}, /* 0x2c9a */
            {8'h00}, /* 0x2c99 */
            {8'h00}, /* 0x2c98 */
            {8'h00}, /* 0x2c97 */
            {8'h00}, /* 0x2c96 */
            {8'h00}, /* 0x2c95 */
            {8'h00}, /* 0x2c94 */
            {8'h00}, /* 0x2c93 */
            {8'h00}, /* 0x2c92 */
            {8'h00}, /* 0x2c91 */
            {8'h00}, /* 0x2c90 */
            {8'h00}, /* 0x2c8f */
            {8'h00}, /* 0x2c8e */
            {8'h00}, /* 0x2c8d */
            {8'h00}, /* 0x2c8c */
            {8'h00}, /* 0x2c8b */
            {8'h00}, /* 0x2c8a */
            {8'h00}, /* 0x2c89 */
            {8'h00}, /* 0x2c88 */
            {8'h00}, /* 0x2c87 */
            {8'h00}, /* 0x2c86 */
            {8'h00}, /* 0x2c85 */
            {8'h00}, /* 0x2c84 */
            {8'h00}, /* 0x2c83 */
            {8'h00}, /* 0x2c82 */
            {8'h00}, /* 0x2c81 */
            {8'h00}, /* 0x2c80 */
            {8'h00}, /* 0x2c7f */
            {8'h00}, /* 0x2c7e */
            {8'h00}, /* 0x2c7d */
            {8'h00}, /* 0x2c7c */
            {8'h00}, /* 0x2c7b */
            {8'h00}, /* 0x2c7a */
            {8'h00}, /* 0x2c79 */
            {8'h00}, /* 0x2c78 */
            {8'h00}, /* 0x2c77 */
            {8'h00}, /* 0x2c76 */
            {8'h00}, /* 0x2c75 */
            {8'h00}, /* 0x2c74 */
            {8'h00}, /* 0x2c73 */
            {8'h00}, /* 0x2c72 */
            {8'h00}, /* 0x2c71 */
            {8'h00}, /* 0x2c70 */
            {8'h00}, /* 0x2c6f */
            {8'h00}, /* 0x2c6e */
            {8'h00}, /* 0x2c6d */
            {8'h00}, /* 0x2c6c */
            {8'h00}, /* 0x2c6b */
            {8'h00}, /* 0x2c6a */
            {8'h00}, /* 0x2c69 */
            {8'h00}, /* 0x2c68 */
            {8'h00}, /* 0x2c67 */
            {8'h00}, /* 0x2c66 */
            {8'h00}, /* 0x2c65 */
            {8'h00}, /* 0x2c64 */
            {8'h00}, /* 0x2c63 */
            {8'h00}, /* 0x2c62 */
            {8'h00}, /* 0x2c61 */
            {8'h00}, /* 0x2c60 */
            {8'h00}, /* 0x2c5f */
            {8'h00}, /* 0x2c5e */
            {8'h00}, /* 0x2c5d */
            {8'h00}, /* 0x2c5c */
            {8'h00}, /* 0x2c5b */
            {8'h00}, /* 0x2c5a */
            {8'h00}, /* 0x2c59 */
            {8'h00}, /* 0x2c58 */
            {8'h00}, /* 0x2c57 */
            {8'h00}, /* 0x2c56 */
            {8'h00}, /* 0x2c55 */
            {8'h00}, /* 0x2c54 */
            {8'h00}, /* 0x2c53 */
            {8'h00}, /* 0x2c52 */
            {8'h00}, /* 0x2c51 */
            {8'h00}, /* 0x2c50 */
            {8'h00}, /* 0x2c4f */
            {8'h00}, /* 0x2c4e */
            {8'h00}, /* 0x2c4d */
            {8'h00}, /* 0x2c4c */
            {8'h00}, /* 0x2c4b */
            {8'h00}, /* 0x2c4a */
            {8'h00}, /* 0x2c49 */
            {8'h00}, /* 0x2c48 */
            {8'h00}, /* 0x2c47 */
            {8'h00}, /* 0x2c46 */
            {8'h00}, /* 0x2c45 */
            {8'h00}, /* 0x2c44 */
            {8'h00}, /* 0x2c43 */
            {8'h00}, /* 0x2c42 */
            {8'h00}, /* 0x2c41 */
            {8'h00}, /* 0x2c40 */
            {8'h00}, /* 0x2c3f */
            {8'h00}, /* 0x2c3e */
            {8'h00}, /* 0x2c3d */
            {8'h00}, /* 0x2c3c */
            {8'h00}, /* 0x2c3b */
            {8'h00}, /* 0x2c3a */
            {8'h00}, /* 0x2c39 */
            {8'h00}, /* 0x2c38 */
            {8'h00}, /* 0x2c37 */
            {8'h00}, /* 0x2c36 */
            {8'h00}, /* 0x2c35 */
            {8'h00}, /* 0x2c34 */
            {8'h00}, /* 0x2c33 */
            {8'h00}, /* 0x2c32 */
            {8'h00}, /* 0x2c31 */
            {8'h00}, /* 0x2c30 */
            {8'h00}, /* 0x2c2f */
            {8'h00}, /* 0x2c2e */
            {8'h00}, /* 0x2c2d */
            {8'h00}, /* 0x2c2c */
            {8'h00}, /* 0x2c2b */
            {8'h00}, /* 0x2c2a */
            {8'h00}, /* 0x2c29 */
            {8'h00}, /* 0x2c28 */
            {8'h00}, /* 0x2c27 */
            {8'h00}, /* 0x2c26 */
            {8'h00}, /* 0x2c25 */
            {8'h00}, /* 0x2c24 */
            {8'h00}, /* 0x2c23 */
            {8'h00}, /* 0x2c22 */
            {8'h00}, /* 0x2c21 */
            {8'h00}, /* 0x2c20 */
            {8'h00}, /* 0x2c1f */
            {8'h00}, /* 0x2c1e */
            {8'h00}, /* 0x2c1d */
            {8'h00}, /* 0x2c1c */
            {8'h00}, /* 0x2c1b */
            {8'h00}, /* 0x2c1a */
            {8'h00}, /* 0x2c19 */
            {8'h00}, /* 0x2c18 */
            {8'h00}, /* 0x2c17 */
            {8'h00}, /* 0x2c16 */
            {8'h00}, /* 0x2c15 */
            {8'h00}, /* 0x2c14 */
            {8'h00}, /* 0x2c13 */
            {8'h00}, /* 0x2c12 */
            {8'h00}, /* 0x2c11 */
            {8'h00}, /* 0x2c10 */
            {8'h00}, /* 0x2c0f */
            {8'h00}, /* 0x2c0e */
            {8'h00}, /* 0x2c0d */
            {8'h00}, /* 0x2c0c */
            {8'h00}, /* 0x2c0b */
            {8'h00}, /* 0x2c0a */
            {8'h00}, /* 0x2c09 */
            {8'h00}, /* 0x2c08 */
            {8'h00}, /* 0x2c07 */
            {8'h00}, /* 0x2c06 */
            {8'h00}, /* 0x2c05 */
            {8'h00}, /* 0x2c04 */
            {8'h00}, /* 0x2c03 */
            {8'h00}, /* 0x2c02 */
            {8'h00}, /* 0x2c01 */
            {8'h00}, /* 0x2c00 */
            {8'h00}, /* 0x2bff */
            {8'h00}, /* 0x2bfe */
            {8'h00}, /* 0x2bfd */
            {8'h00}, /* 0x2bfc */
            {8'h00}, /* 0x2bfb */
            {8'h00}, /* 0x2bfa */
            {8'h00}, /* 0x2bf9 */
            {8'h00}, /* 0x2bf8 */
            {8'h00}, /* 0x2bf7 */
            {8'h00}, /* 0x2bf6 */
            {8'h00}, /* 0x2bf5 */
            {8'h00}, /* 0x2bf4 */
            {8'h00}, /* 0x2bf3 */
            {8'h00}, /* 0x2bf2 */
            {8'h00}, /* 0x2bf1 */
            {8'h00}, /* 0x2bf0 */
            {8'h00}, /* 0x2bef */
            {8'h00}, /* 0x2bee */
            {8'h00}, /* 0x2bed */
            {8'h00}, /* 0x2bec */
            {8'h00}, /* 0x2beb */
            {8'h00}, /* 0x2bea */
            {8'h00}, /* 0x2be9 */
            {8'h00}, /* 0x2be8 */
            {8'h00}, /* 0x2be7 */
            {8'h00}, /* 0x2be6 */
            {8'h00}, /* 0x2be5 */
            {8'h00}, /* 0x2be4 */
            {8'h00}, /* 0x2be3 */
            {8'h00}, /* 0x2be2 */
            {8'h00}, /* 0x2be1 */
            {8'h00}, /* 0x2be0 */
            {8'h00}, /* 0x2bdf */
            {8'h00}, /* 0x2bde */
            {8'h00}, /* 0x2bdd */
            {8'h00}, /* 0x2bdc */
            {8'h00}, /* 0x2bdb */
            {8'h00}, /* 0x2bda */
            {8'h00}, /* 0x2bd9 */
            {8'h00}, /* 0x2bd8 */
            {8'h00}, /* 0x2bd7 */
            {8'h00}, /* 0x2bd6 */
            {8'h00}, /* 0x2bd5 */
            {8'h00}, /* 0x2bd4 */
            {8'h00}, /* 0x2bd3 */
            {8'h00}, /* 0x2bd2 */
            {8'h00}, /* 0x2bd1 */
            {8'h00}, /* 0x2bd0 */
            {8'h00}, /* 0x2bcf */
            {8'h00}, /* 0x2bce */
            {8'h00}, /* 0x2bcd */
            {8'h00}, /* 0x2bcc */
            {8'h00}, /* 0x2bcb */
            {8'h00}, /* 0x2bca */
            {8'h00}, /* 0x2bc9 */
            {8'h00}, /* 0x2bc8 */
            {8'h00}, /* 0x2bc7 */
            {8'h00}, /* 0x2bc6 */
            {8'h00}, /* 0x2bc5 */
            {8'h00}, /* 0x2bc4 */
            {8'h00}, /* 0x2bc3 */
            {8'h00}, /* 0x2bc2 */
            {8'h00}, /* 0x2bc1 */
            {8'h00}, /* 0x2bc0 */
            {8'h00}, /* 0x2bbf */
            {8'h00}, /* 0x2bbe */
            {8'h00}, /* 0x2bbd */
            {8'h00}, /* 0x2bbc */
            {8'h00}, /* 0x2bbb */
            {8'h00}, /* 0x2bba */
            {8'h00}, /* 0x2bb9 */
            {8'h00}, /* 0x2bb8 */
            {8'h00}, /* 0x2bb7 */
            {8'h00}, /* 0x2bb6 */
            {8'h00}, /* 0x2bb5 */
            {8'h00}, /* 0x2bb4 */
            {8'h00}, /* 0x2bb3 */
            {8'h00}, /* 0x2bb2 */
            {8'h00}, /* 0x2bb1 */
            {8'h00}, /* 0x2bb0 */
            {8'h00}, /* 0x2baf */
            {8'h00}, /* 0x2bae */
            {8'h00}, /* 0x2bad */
            {8'h00}, /* 0x2bac */
            {8'h00}, /* 0x2bab */
            {8'h00}, /* 0x2baa */
            {8'h00}, /* 0x2ba9 */
            {8'h00}, /* 0x2ba8 */
            {8'h00}, /* 0x2ba7 */
            {8'h00}, /* 0x2ba6 */
            {8'h00}, /* 0x2ba5 */
            {8'h00}, /* 0x2ba4 */
            {8'h00}, /* 0x2ba3 */
            {8'h00}, /* 0x2ba2 */
            {8'h00}, /* 0x2ba1 */
            {8'h00}, /* 0x2ba0 */
            {8'h00}, /* 0x2b9f */
            {8'h00}, /* 0x2b9e */
            {8'h00}, /* 0x2b9d */
            {8'h00}, /* 0x2b9c */
            {8'h00}, /* 0x2b9b */
            {8'h00}, /* 0x2b9a */
            {8'h00}, /* 0x2b99 */
            {8'h00}, /* 0x2b98 */
            {8'h00}, /* 0x2b97 */
            {8'h00}, /* 0x2b96 */
            {8'h00}, /* 0x2b95 */
            {8'h00}, /* 0x2b94 */
            {8'h00}, /* 0x2b93 */
            {8'h00}, /* 0x2b92 */
            {8'h00}, /* 0x2b91 */
            {8'h00}, /* 0x2b90 */
            {8'h00}, /* 0x2b8f */
            {8'h00}, /* 0x2b8e */
            {8'h00}, /* 0x2b8d */
            {8'h00}, /* 0x2b8c */
            {8'h00}, /* 0x2b8b */
            {8'h00}, /* 0x2b8a */
            {8'h00}, /* 0x2b89 */
            {8'h00}, /* 0x2b88 */
            {8'h00}, /* 0x2b87 */
            {8'h00}, /* 0x2b86 */
            {8'h00}, /* 0x2b85 */
            {8'h00}, /* 0x2b84 */
            {8'h00}, /* 0x2b83 */
            {8'h00}, /* 0x2b82 */
            {8'h00}, /* 0x2b81 */
            {8'h00}, /* 0x2b80 */
            {8'h00}, /* 0x2b7f */
            {8'h00}, /* 0x2b7e */
            {8'h00}, /* 0x2b7d */
            {8'h00}, /* 0x2b7c */
            {8'h00}, /* 0x2b7b */
            {8'h00}, /* 0x2b7a */
            {8'h00}, /* 0x2b79 */
            {8'h00}, /* 0x2b78 */
            {8'h00}, /* 0x2b77 */
            {8'h00}, /* 0x2b76 */
            {8'h00}, /* 0x2b75 */
            {8'h00}, /* 0x2b74 */
            {8'h00}, /* 0x2b73 */
            {8'h00}, /* 0x2b72 */
            {8'h00}, /* 0x2b71 */
            {8'h00}, /* 0x2b70 */
            {8'h00}, /* 0x2b6f */
            {8'h00}, /* 0x2b6e */
            {8'h00}, /* 0x2b6d */
            {8'h00}, /* 0x2b6c */
            {8'h00}, /* 0x2b6b */
            {8'h00}, /* 0x2b6a */
            {8'h00}, /* 0x2b69 */
            {8'h00}, /* 0x2b68 */
            {8'h00}, /* 0x2b67 */
            {8'h00}, /* 0x2b66 */
            {8'h00}, /* 0x2b65 */
            {8'h00}, /* 0x2b64 */
            {8'h00}, /* 0x2b63 */
            {8'h00}, /* 0x2b62 */
            {8'h00}, /* 0x2b61 */
            {8'h00}, /* 0x2b60 */
            {8'h00}, /* 0x2b5f */
            {8'h00}, /* 0x2b5e */
            {8'h00}, /* 0x2b5d */
            {8'h00}, /* 0x2b5c */
            {8'h00}, /* 0x2b5b */
            {8'h00}, /* 0x2b5a */
            {8'h00}, /* 0x2b59 */
            {8'h00}, /* 0x2b58 */
            {8'h00}, /* 0x2b57 */
            {8'h00}, /* 0x2b56 */
            {8'h00}, /* 0x2b55 */
            {8'h00}, /* 0x2b54 */
            {8'h00}, /* 0x2b53 */
            {8'h00}, /* 0x2b52 */
            {8'h00}, /* 0x2b51 */
            {8'h00}, /* 0x2b50 */
            {8'h00}, /* 0x2b4f */
            {8'h00}, /* 0x2b4e */
            {8'h00}, /* 0x2b4d */
            {8'h00}, /* 0x2b4c */
            {8'h00}, /* 0x2b4b */
            {8'h00}, /* 0x2b4a */
            {8'h00}, /* 0x2b49 */
            {8'h00}, /* 0x2b48 */
            {8'h00}, /* 0x2b47 */
            {8'h00}, /* 0x2b46 */
            {8'h00}, /* 0x2b45 */
            {8'h00}, /* 0x2b44 */
            {8'h00}, /* 0x2b43 */
            {8'h00}, /* 0x2b42 */
            {8'h00}, /* 0x2b41 */
            {8'h00}, /* 0x2b40 */
            {8'h00}, /* 0x2b3f */
            {8'h00}, /* 0x2b3e */
            {8'h00}, /* 0x2b3d */
            {8'h00}, /* 0x2b3c */
            {8'h00}, /* 0x2b3b */
            {8'h00}, /* 0x2b3a */
            {8'h00}, /* 0x2b39 */
            {8'h00}, /* 0x2b38 */
            {8'h00}, /* 0x2b37 */
            {8'h00}, /* 0x2b36 */
            {8'h00}, /* 0x2b35 */
            {8'h00}, /* 0x2b34 */
            {8'h00}, /* 0x2b33 */
            {8'h00}, /* 0x2b32 */
            {8'h00}, /* 0x2b31 */
            {8'h00}, /* 0x2b30 */
            {8'h00}, /* 0x2b2f */
            {8'h00}, /* 0x2b2e */
            {8'h00}, /* 0x2b2d */
            {8'h00}, /* 0x2b2c */
            {8'h00}, /* 0x2b2b */
            {8'h00}, /* 0x2b2a */
            {8'h00}, /* 0x2b29 */
            {8'h00}, /* 0x2b28 */
            {8'h00}, /* 0x2b27 */
            {8'h00}, /* 0x2b26 */
            {8'h00}, /* 0x2b25 */
            {8'h00}, /* 0x2b24 */
            {8'h00}, /* 0x2b23 */
            {8'h00}, /* 0x2b22 */
            {8'h00}, /* 0x2b21 */
            {8'h00}, /* 0x2b20 */
            {8'h00}, /* 0x2b1f */
            {8'h00}, /* 0x2b1e */
            {8'h00}, /* 0x2b1d */
            {8'h00}, /* 0x2b1c */
            {8'h00}, /* 0x2b1b */
            {8'h00}, /* 0x2b1a */
            {8'h00}, /* 0x2b19 */
            {8'h00}, /* 0x2b18 */
            {8'h00}, /* 0x2b17 */
            {8'h00}, /* 0x2b16 */
            {8'h00}, /* 0x2b15 */
            {8'h00}, /* 0x2b14 */
            {8'h00}, /* 0x2b13 */
            {8'h00}, /* 0x2b12 */
            {8'h00}, /* 0x2b11 */
            {8'h00}, /* 0x2b10 */
            {8'h00}, /* 0x2b0f */
            {8'h00}, /* 0x2b0e */
            {8'h00}, /* 0x2b0d */
            {8'h00}, /* 0x2b0c */
            {8'h00}, /* 0x2b0b */
            {8'h00}, /* 0x2b0a */
            {8'h00}, /* 0x2b09 */
            {8'h00}, /* 0x2b08 */
            {8'h00}, /* 0x2b07 */
            {8'h00}, /* 0x2b06 */
            {8'h00}, /* 0x2b05 */
            {8'h00}, /* 0x2b04 */
            {8'h00}, /* 0x2b03 */
            {8'h00}, /* 0x2b02 */
            {8'h00}, /* 0x2b01 */
            {8'h00}, /* 0x2b00 */
            {8'h00}, /* 0x2aff */
            {8'h00}, /* 0x2afe */
            {8'h00}, /* 0x2afd */
            {8'h00}, /* 0x2afc */
            {8'h00}, /* 0x2afb */
            {8'h00}, /* 0x2afa */
            {8'h00}, /* 0x2af9 */
            {8'h00}, /* 0x2af8 */
            {8'h00}, /* 0x2af7 */
            {8'h00}, /* 0x2af6 */
            {8'h00}, /* 0x2af5 */
            {8'h00}, /* 0x2af4 */
            {8'h00}, /* 0x2af3 */
            {8'h00}, /* 0x2af2 */
            {8'h00}, /* 0x2af1 */
            {8'h00}, /* 0x2af0 */
            {8'h00}, /* 0x2aef */
            {8'h00}, /* 0x2aee */
            {8'h00}, /* 0x2aed */
            {8'h00}, /* 0x2aec */
            {8'h00}, /* 0x2aeb */
            {8'h00}, /* 0x2aea */
            {8'h00}, /* 0x2ae9 */
            {8'h00}, /* 0x2ae8 */
            {8'h00}, /* 0x2ae7 */
            {8'h00}, /* 0x2ae6 */
            {8'h00}, /* 0x2ae5 */
            {8'h00}, /* 0x2ae4 */
            {8'h00}, /* 0x2ae3 */
            {8'h00}, /* 0x2ae2 */
            {8'h00}, /* 0x2ae1 */
            {8'h00}, /* 0x2ae0 */
            {8'h00}, /* 0x2adf */
            {8'h00}, /* 0x2ade */
            {8'h00}, /* 0x2add */
            {8'h00}, /* 0x2adc */
            {8'h00}, /* 0x2adb */
            {8'h00}, /* 0x2ada */
            {8'h00}, /* 0x2ad9 */
            {8'h00}, /* 0x2ad8 */
            {8'h00}, /* 0x2ad7 */
            {8'h00}, /* 0x2ad6 */
            {8'h00}, /* 0x2ad5 */
            {8'h00}, /* 0x2ad4 */
            {8'h00}, /* 0x2ad3 */
            {8'h00}, /* 0x2ad2 */
            {8'h00}, /* 0x2ad1 */
            {8'h00}, /* 0x2ad0 */
            {8'h00}, /* 0x2acf */
            {8'h00}, /* 0x2ace */
            {8'h00}, /* 0x2acd */
            {8'h00}, /* 0x2acc */
            {8'h00}, /* 0x2acb */
            {8'h00}, /* 0x2aca */
            {8'h00}, /* 0x2ac9 */
            {8'h00}, /* 0x2ac8 */
            {8'h00}, /* 0x2ac7 */
            {8'h00}, /* 0x2ac6 */
            {8'h00}, /* 0x2ac5 */
            {8'h00}, /* 0x2ac4 */
            {8'h00}, /* 0x2ac3 */
            {8'h00}, /* 0x2ac2 */
            {8'h00}, /* 0x2ac1 */
            {8'h00}, /* 0x2ac0 */
            {8'h00}, /* 0x2abf */
            {8'h00}, /* 0x2abe */
            {8'h00}, /* 0x2abd */
            {8'h00}, /* 0x2abc */
            {8'h00}, /* 0x2abb */
            {8'h00}, /* 0x2aba */
            {8'h00}, /* 0x2ab9 */
            {8'h00}, /* 0x2ab8 */
            {8'h00}, /* 0x2ab7 */
            {8'h00}, /* 0x2ab6 */
            {8'h00}, /* 0x2ab5 */
            {8'h00}, /* 0x2ab4 */
            {8'h00}, /* 0x2ab3 */
            {8'h00}, /* 0x2ab2 */
            {8'h00}, /* 0x2ab1 */
            {8'h00}, /* 0x2ab0 */
            {8'h00}, /* 0x2aaf */
            {8'h00}, /* 0x2aae */
            {8'h00}, /* 0x2aad */
            {8'h00}, /* 0x2aac */
            {8'h00}, /* 0x2aab */
            {8'h00}, /* 0x2aaa */
            {8'h00}, /* 0x2aa9 */
            {8'h00}, /* 0x2aa8 */
            {8'h00}, /* 0x2aa7 */
            {8'h00}, /* 0x2aa6 */
            {8'h00}, /* 0x2aa5 */
            {8'h00}, /* 0x2aa4 */
            {8'h00}, /* 0x2aa3 */
            {8'h00}, /* 0x2aa2 */
            {8'h00}, /* 0x2aa1 */
            {8'h00}, /* 0x2aa0 */
            {8'h00}, /* 0x2a9f */
            {8'h00}, /* 0x2a9e */
            {8'h00}, /* 0x2a9d */
            {8'h00}, /* 0x2a9c */
            {8'h00}, /* 0x2a9b */
            {8'h00}, /* 0x2a9a */
            {8'h00}, /* 0x2a99 */
            {8'h00}, /* 0x2a98 */
            {8'h00}, /* 0x2a97 */
            {8'h00}, /* 0x2a96 */
            {8'h00}, /* 0x2a95 */
            {8'h00}, /* 0x2a94 */
            {8'h00}, /* 0x2a93 */
            {8'h00}, /* 0x2a92 */
            {8'h00}, /* 0x2a91 */
            {8'h00}, /* 0x2a90 */
            {8'h00}, /* 0x2a8f */
            {8'h00}, /* 0x2a8e */
            {8'h00}, /* 0x2a8d */
            {8'h00}, /* 0x2a8c */
            {8'h00}, /* 0x2a8b */
            {8'h00}, /* 0x2a8a */
            {8'h00}, /* 0x2a89 */
            {8'h00}, /* 0x2a88 */
            {8'h00}, /* 0x2a87 */
            {8'h00}, /* 0x2a86 */
            {8'h00}, /* 0x2a85 */
            {8'h00}, /* 0x2a84 */
            {8'h00}, /* 0x2a83 */
            {8'h00}, /* 0x2a82 */
            {8'h00}, /* 0x2a81 */
            {8'h00}, /* 0x2a80 */
            {8'h00}, /* 0x2a7f */
            {8'h00}, /* 0x2a7e */
            {8'h00}, /* 0x2a7d */
            {8'h00}, /* 0x2a7c */
            {8'h00}, /* 0x2a7b */
            {8'h00}, /* 0x2a7a */
            {8'h00}, /* 0x2a79 */
            {8'h00}, /* 0x2a78 */
            {8'h00}, /* 0x2a77 */
            {8'h00}, /* 0x2a76 */
            {8'h00}, /* 0x2a75 */
            {8'h00}, /* 0x2a74 */
            {8'h00}, /* 0x2a73 */
            {8'h00}, /* 0x2a72 */
            {8'h00}, /* 0x2a71 */
            {8'h00}, /* 0x2a70 */
            {8'h00}, /* 0x2a6f */
            {8'h00}, /* 0x2a6e */
            {8'h00}, /* 0x2a6d */
            {8'h00}, /* 0x2a6c */
            {8'h00}, /* 0x2a6b */
            {8'h00}, /* 0x2a6a */
            {8'h00}, /* 0x2a69 */
            {8'h00}, /* 0x2a68 */
            {8'h00}, /* 0x2a67 */
            {8'h00}, /* 0x2a66 */
            {8'h00}, /* 0x2a65 */
            {8'h00}, /* 0x2a64 */
            {8'h00}, /* 0x2a63 */
            {8'h00}, /* 0x2a62 */
            {8'h00}, /* 0x2a61 */
            {8'h00}, /* 0x2a60 */
            {8'h00}, /* 0x2a5f */
            {8'h00}, /* 0x2a5e */
            {8'h00}, /* 0x2a5d */
            {8'h00}, /* 0x2a5c */
            {8'h00}, /* 0x2a5b */
            {8'h00}, /* 0x2a5a */
            {8'h00}, /* 0x2a59 */
            {8'h00}, /* 0x2a58 */
            {8'h00}, /* 0x2a57 */
            {8'h00}, /* 0x2a56 */
            {8'h00}, /* 0x2a55 */
            {8'h00}, /* 0x2a54 */
            {8'h00}, /* 0x2a53 */
            {8'h00}, /* 0x2a52 */
            {8'h00}, /* 0x2a51 */
            {8'h00}, /* 0x2a50 */
            {8'h00}, /* 0x2a4f */
            {8'h00}, /* 0x2a4e */
            {8'h00}, /* 0x2a4d */
            {8'h00}, /* 0x2a4c */
            {8'h00}, /* 0x2a4b */
            {8'h00}, /* 0x2a4a */
            {8'h00}, /* 0x2a49 */
            {8'h00}, /* 0x2a48 */
            {8'h00}, /* 0x2a47 */
            {8'h00}, /* 0x2a46 */
            {8'h00}, /* 0x2a45 */
            {8'h00}, /* 0x2a44 */
            {8'h00}, /* 0x2a43 */
            {8'h00}, /* 0x2a42 */
            {8'h00}, /* 0x2a41 */
            {8'h00}, /* 0x2a40 */
            {8'h00}, /* 0x2a3f */
            {8'h00}, /* 0x2a3e */
            {8'h00}, /* 0x2a3d */
            {8'h00}, /* 0x2a3c */
            {8'h00}, /* 0x2a3b */
            {8'h00}, /* 0x2a3a */
            {8'h00}, /* 0x2a39 */
            {8'h00}, /* 0x2a38 */
            {8'h00}, /* 0x2a37 */
            {8'h00}, /* 0x2a36 */
            {8'h00}, /* 0x2a35 */
            {8'h00}, /* 0x2a34 */
            {8'h00}, /* 0x2a33 */
            {8'h00}, /* 0x2a32 */
            {8'h00}, /* 0x2a31 */
            {8'h00}, /* 0x2a30 */
            {8'h00}, /* 0x2a2f */
            {8'h00}, /* 0x2a2e */
            {8'h00}, /* 0x2a2d */
            {8'h00}, /* 0x2a2c */
            {8'h00}, /* 0x2a2b */
            {8'h00}, /* 0x2a2a */
            {8'h00}, /* 0x2a29 */
            {8'h00}, /* 0x2a28 */
            {8'h00}, /* 0x2a27 */
            {8'h00}, /* 0x2a26 */
            {8'h00}, /* 0x2a25 */
            {8'h00}, /* 0x2a24 */
            {8'h00}, /* 0x2a23 */
            {8'h00}, /* 0x2a22 */
            {8'h00}, /* 0x2a21 */
            {8'h00}, /* 0x2a20 */
            {8'h00}, /* 0x2a1f */
            {8'h00}, /* 0x2a1e */
            {8'h00}, /* 0x2a1d */
            {8'h00}, /* 0x2a1c */
            {8'h00}, /* 0x2a1b */
            {8'h00}, /* 0x2a1a */
            {8'h00}, /* 0x2a19 */
            {8'h00}, /* 0x2a18 */
            {8'h00}, /* 0x2a17 */
            {8'h00}, /* 0x2a16 */
            {8'h00}, /* 0x2a15 */
            {8'h00}, /* 0x2a14 */
            {8'h00}, /* 0x2a13 */
            {8'h00}, /* 0x2a12 */
            {8'h00}, /* 0x2a11 */
            {8'h00}, /* 0x2a10 */
            {8'h00}, /* 0x2a0f */
            {8'h00}, /* 0x2a0e */
            {8'h00}, /* 0x2a0d */
            {8'h00}, /* 0x2a0c */
            {8'h00}, /* 0x2a0b */
            {8'h00}, /* 0x2a0a */
            {8'h00}, /* 0x2a09 */
            {8'h00}, /* 0x2a08 */
            {8'h00}, /* 0x2a07 */
            {8'h00}, /* 0x2a06 */
            {8'h00}, /* 0x2a05 */
            {8'h00}, /* 0x2a04 */
            {8'h00}, /* 0x2a03 */
            {8'h00}, /* 0x2a02 */
            {8'h00}, /* 0x2a01 */
            {8'h00}, /* 0x2a00 */
            {8'h00}, /* 0x29ff */
            {8'h00}, /* 0x29fe */
            {8'h00}, /* 0x29fd */
            {8'h00}, /* 0x29fc */
            {8'h00}, /* 0x29fb */
            {8'h00}, /* 0x29fa */
            {8'h00}, /* 0x29f9 */
            {8'h00}, /* 0x29f8 */
            {8'h00}, /* 0x29f7 */
            {8'h00}, /* 0x29f6 */
            {8'h00}, /* 0x29f5 */
            {8'h00}, /* 0x29f4 */
            {8'h00}, /* 0x29f3 */
            {8'h00}, /* 0x29f2 */
            {8'h00}, /* 0x29f1 */
            {8'h00}, /* 0x29f0 */
            {8'h00}, /* 0x29ef */
            {8'h00}, /* 0x29ee */
            {8'h00}, /* 0x29ed */
            {8'h00}, /* 0x29ec */
            {8'h00}, /* 0x29eb */
            {8'h00}, /* 0x29ea */
            {8'h00}, /* 0x29e9 */
            {8'h00}, /* 0x29e8 */
            {8'h00}, /* 0x29e7 */
            {8'h00}, /* 0x29e6 */
            {8'h00}, /* 0x29e5 */
            {8'h00}, /* 0x29e4 */
            {8'h00}, /* 0x29e3 */
            {8'h00}, /* 0x29e2 */
            {8'h00}, /* 0x29e1 */
            {8'h00}, /* 0x29e0 */
            {8'h00}, /* 0x29df */
            {8'h00}, /* 0x29de */
            {8'h00}, /* 0x29dd */
            {8'h00}, /* 0x29dc */
            {8'h00}, /* 0x29db */
            {8'h00}, /* 0x29da */
            {8'h00}, /* 0x29d9 */
            {8'h00}, /* 0x29d8 */
            {8'h00}, /* 0x29d7 */
            {8'h00}, /* 0x29d6 */
            {8'h00}, /* 0x29d5 */
            {8'h00}, /* 0x29d4 */
            {8'h00}, /* 0x29d3 */
            {8'h00}, /* 0x29d2 */
            {8'h00}, /* 0x29d1 */
            {8'h00}, /* 0x29d0 */
            {8'h00}, /* 0x29cf */
            {8'h00}, /* 0x29ce */
            {8'h00}, /* 0x29cd */
            {8'h00}, /* 0x29cc */
            {8'h00}, /* 0x29cb */
            {8'h00}, /* 0x29ca */
            {8'h00}, /* 0x29c9 */
            {8'h00}, /* 0x29c8 */
            {8'h00}, /* 0x29c7 */
            {8'h00}, /* 0x29c6 */
            {8'h00}, /* 0x29c5 */
            {8'h00}, /* 0x29c4 */
            {8'h00}, /* 0x29c3 */
            {8'h00}, /* 0x29c2 */
            {8'h00}, /* 0x29c1 */
            {8'h00}, /* 0x29c0 */
            {8'h00}, /* 0x29bf */
            {8'h00}, /* 0x29be */
            {8'h00}, /* 0x29bd */
            {8'h00}, /* 0x29bc */
            {8'h00}, /* 0x29bb */
            {8'h00}, /* 0x29ba */
            {8'h00}, /* 0x29b9 */
            {8'h00}, /* 0x29b8 */
            {8'h00}, /* 0x29b7 */
            {8'h00}, /* 0x29b6 */
            {8'h00}, /* 0x29b5 */
            {8'h00}, /* 0x29b4 */
            {8'h00}, /* 0x29b3 */
            {8'h00}, /* 0x29b2 */
            {8'h00}, /* 0x29b1 */
            {8'h00}, /* 0x29b0 */
            {8'h00}, /* 0x29af */
            {8'h00}, /* 0x29ae */
            {8'h00}, /* 0x29ad */
            {8'h00}, /* 0x29ac */
            {8'h00}, /* 0x29ab */
            {8'h00}, /* 0x29aa */
            {8'h00}, /* 0x29a9 */
            {8'h00}, /* 0x29a8 */
            {8'h00}, /* 0x29a7 */
            {8'h00}, /* 0x29a6 */
            {8'h00}, /* 0x29a5 */
            {8'h00}, /* 0x29a4 */
            {8'h00}, /* 0x29a3 */
            {8'h00}, /* 0x29a2 */
            {8'h00}, /* 0x29a1 */
            {8'h00}, /* 0x29a0 */
            {8'h00}, /* 0x299f */
            {8'h00}, /* 0x299e */
            {8'h00}, /* 0x299d */
            {8'h00}, /* 0x299c */
            {8'h00}, /* 0x299b */
            {8'h00}, /* 0x299a */
            {8'h00}, /* 0x2999 */
            {8'h00}, /* 0x2998 */
            {8'h00}, /* 0x2997 */
            {8'h00}, /* 0x2996 */
            {8'h00}, /* 0x2995 */
            {8'h00}, /* 0x2994 */
            {8'h00}, /* 0x2993 */
            {8'h00}, /* 0x2992 */
            {8'h00}, /* 0x2991 */
            {8'h00}, /* 0x2990 */
            {8'h00}, /* 0x298f */
            {8'h00}, /* 0x298e */
            {8'h00}, /* 0x298d */
            {8'h00}, /* 0x298c */
            {8'h00}, /* 0x298b */
            {8'h00}, /* 0x298a */
            {8'h00}, /* 0x2989 */
            {8'h00}, /* 0x2988 */
            {8'h00}, /* 0x2987 */
            {8'h00}, /* 0x2986 */
            {8'h00}, /* 0x2985 */
            {8'h00}, /* 0x2984 */
            {8'h00}, /* 0x2983 */
            {8'h00}, /* 0x2982 */
            {8'h00}, /* 0x2981 */
            {8'h00}, /* 0x2980 */
            {8'h00}, /* 0x297f */
            {8'h00}, /* 0x297e */
            {8'h00}, /* 0x297d */
            {8'h00}, /* 0x297c */
            {8'h00}, /* 0x297b */
            {8'h00}, /* 0x297a */
            {8'h00}, /* 0x2979 */
            {8'h00}, /* 0x2978 */
            {8'h00}, /* 0x2977 */
            {8'h00}, /* 0x2976 */
            {8'h00}, /* 0x2975 */
            {8'h00}, /* 0x2974 */
            {8'h00}, /* 0x2973 */
            {8'h00}, /* 0x2972 */
            {8'h00}, /* 0x2971 */
            {8'h00}, /* 0x2970 */
            {8'h00}, /* 0x296f */
            {8'h00}, /* 0x296e */
            {8'h00}, /* 0x296d */
            {8'h00}, /* 0x296c */
            {8'h00}, /* 0x296b */
            {8'h00}, /* 0x296a */
            {8'h00}, /* 0x2969 */
            {8'h00}, /* 0x2968 */
            {8'h00}, /* 0x2967 */
            {8'h00}, /* 0x2966 */
            {8'h00}, /* 0x2965 */
            {8'h00}, /* 0x2964 */
            {8'h00}, /* 0x2963 */
            {8'h00}, /* 0x2962 */
            {8'h00}, /* 0x2961 */
            {8'h00}, /* 0x2960 */
            {8'h00}, /* 0x295f */
            {8'h00}, /* 0x295e */
            {8'h00}, /* 0x295d */
            {8'h00}, /* 0x295c */
            {8'h00}, /* 0x295b */
            {8'h00}, /* 0x295a */
            {8'h00}, /* 0x2959 */
            {8'h00}, /* 0x2958 */
            {8'h00}, /* 0x2957 */
            {8'h00}, /* 0x2956 */
            {8'h00}, /* 0x2955 */
            {8'h00}, /* 0x2954 */
            {8'h00}, /* 0x2953 */
            {8'h00}, /* 0x2952 */
            {8'h00}, /* 0x2951 */
            {8'h00}, /* 0x2950 */
            {8'h00}, /* 0x294f */
            {8'h00}, /* 0x294e */
            {8'h00}, /* 0x294d */
            {8'h00}, /* 0x294c */
            {8'h00}, /* 0x294b */
            {8'h00}, /* 0x294a */
            {8'h00}, /* 0x2949 */
            {8'h00}, /* 0x2948 */
            {8'h00}, /* 0x2947 */
            {8'h00}, /* 0x2946 */
            {8'h00}, /* 0x2945 */
            {8'h00}, /* 0x2944 */
            {8'h00}, /* 0x2943 */
            {8'h00}, /* 0x2942 */
            {8'h00}, /* 0x2941 */
            {8'h00}, /* 0x2940 */
            {8'h00}, /* 0x293f */
            {8'h00}, /* 0x293e */
            {8'h00}, /* 0x293d */
            {8'h00}, /* 0x293c */
            {8'h00}, /* 0x293b */
            {8'h00}, /* 0x293a */
            {8'h00}, /* 0x2939 */
            {8'h00}, /* 0x2938 */
            {8'h00}, /* 0x2937 */
            {8'h00}, /* 0x2936 */
            {8'h00}, /* 0x2935 */
            {8'h00}, /* 0x2934 */
            {8'h00}, /* 0x2933 */
            {8'h00}, /* 0x2932 */
            {8'h00}, /* 0x2931 */
            {8'h00}, /* 0x2930 */
            {8'h00}, /* 0x292f */
            {8'h00}, /* 0x292e */
            {8'h00}, /* 0x292d */
            {8'h00}, /* 0x292c */
            {8'h00}, /* 0x292b */
            {8'h00}, /* 0x292a */
            {8'h00}, /* 0x2929 */
            {8'h00}, /* 0x2928 */
            {8'h00}, /* 0x2927 */
            {8'h00}, /* 0x2926 */
            {8'h00}, /* 0x2925 */
            {8'h00}, /* 0x2924 */
            {8'h00}, /* 0x2923 */
            {8'h00}, /* 0x2922 */
            {8'h00}, /* 0x2921 */
            {8'h00}, /* 0x2920 */
            {8'h00}, /* 0x291f */
            {8'h00}, /* 0x291e */
            {8'h00}, /* 0x291d */
            {8'h00}, /* 0x291c */
            {8'h00}, /* 0x291b */
            {8'h00}, /* 0x291a */
            {8'h00}, /* 0x2919 */
            {8'h00}, /* 0x2918 */
            {8'h00}, /* 0x2917 */
            {8'h00}, /* 0x2916 */
            {8'h00}, /* 0x2915 */
            {8'h00}, /* 0x2914 */
            {8'h00}, /* 0x2913 */
            {8'h00}, /* 0x2912 */
            {8'h00}, /* 0x2911 */
            {8'h00}, /* 0x2910 */
            {8'h00}, /* 0x290f */
            {8'h00}, /* 0x290e */
            {8'h00}, /* 0x290d */
            {8'h00}, /* 0x290c */
            {8'h00}, /* 0x290b */
            {8'h00}, /* 0x290a */
            {8'h00}, /* 0x2909 */
            {8'h00}, /* 0x2908 */
            {8'h00}, /* 0x2907 */
            {8'h00}, /* 0x2906 */
            {8'h00}, /* 0x2905 */
            {8'h00}, /* 0x2904 */
            {8'h00}, /* 0x2903 */
            {8'h00}, /* 0x2902 */
            {8'h00}, /* 0x2901 */
            {8'h00}, /* 0x2900 */
            {8'h00}, /* 0x28ff */
            {8'h00}, /* 0x28fe */
            {8'h00}, /* 0x28fd */
            {8'h00}, /* 0x28fc */
            {8'h00}, /* 0x28fb */
            {8'h00}, /* 0x28fa */
            {8'h00}, /* 0x28f9 */
            {8'h00}, /* 0x28f8 */
            {8'h00}, /* 0x28f7 */
            {8'h00}, /* 0x28f6 */
            {8'h00}, /* 0x28f5 */
            {8'h00}, /* 0x28f4 */
            {8'h00}, /* 0x28f3 */
            {8'h00}, /* 0x28f2 */
            {8'h00}, /* 0x28f1 */
            {8'h00}, /* 0x28f0 */
            {8'h00}, /* 0x28ef */
            {8'h00}, /* 0x28ee */
            {8'h00}, /* 0x28ed */
            {8'h00}, /* 0x28ec */
            {8'h00}, /* 0x28eb */
            {8'h00}, /* 0x28ea */
            {8'h00}, /* 0x28e9 */
            {8'h00}, /* 0x28e8 */
            {8'h00}, /* 0x28e7 */
            {8'h00}, /* 0x28e6 */
            {8'h00}, /* 0x28e5 */
            {8'h00}, /* 0x28e4 */
            {8'h00}, /* 0x28e3 */
            {8'h00}, /* 0x28e2 */
            {8'h00}, /* 0x28e1 */
            {8'h00}, /* 0x28e0 */
            {8'h00}, /* 0x28df */
            {8'h00}, /* 0x28de */
            {8'h00}, /* 0x28dd */
            {8'h00}, /* 0x28dc */
            {8'h00}, /* 0x28db */
            {8'h00}, /* 0x28da */
            {8'h00}, /* 0x28d9 */
            {8'h00}, /* 0x28d8 */
            {8'h00}, /* 0x28d7 */
            {8'h00}, /* 0x28d6 */
            {8'h00}, /* 0x28d5 */
            {8'h00}, /* 0x28d4 */
            {8'h00}, /* 0x28d3 */
            {8'h00}, /* 0x28d2 */
            {8'h00}, /* 0x28d1 */
            {8'h00}, /* 0x28d0 */
            {8'h00}, /* 0x28cf */
            {8'h00}, /* 0x28ce */
            {8'h00}, /* 0x28cd */
            {8'h00}, /* 0x28cc */
            {8'h00}, /* 0x28cb */
            {8'h00}, /* 0x28ca */
            {8'h00}, /* 0x28c9 */
            {8'h00}, /* 0x28c8 */
            {8'h00}, /* 0x28c7 */
            {8'h00}, /* 0x28c6 */
            {8'h00}, /* 0x28c5 */
            {8'h00}, /* 0x28c4 */
            {8'h00}, /* 0x28c3 */
            {8'h00}, /* 0x28c2 */
            {8'h00}, /* 0x28c1 */
            {8'h00}, /* 0x28c0 */
            {8'h00}, /* 0x28bf */
            {8'h00}, /* 0x28be */
            {8'h00}, /* 0x28bd */
            {8'h00}, /* 0x28bc */
            {8'h00}, /* 0x28bb */
            {8'h00}, /* 0x28ba */
            {8'h00}, /* 0x28b9 */
            {8'h00}, /* 0x28b8 */
            {8'h00}, /* 0x28b7 */
            {8'h00}, /* 0x28b6 */
            {8'h00}, /* 0x28b5 */
            {8'h00}, /* 0x28b4 */
            {8'h00}, /* 0x28b3 */
            {8'h00}, /* 0x28b2 */
            {8'h00}, /* 0x28b1 */
            {8'h00}, /* 0x28b0 */
            {8'h00}, /* 0x28af */
            {8'h00}, /* 0x28ae */
            {8'h00}, /* 0x28ad */
            {8'h00}, /* 0x28ac */
            {8'h00}, /* 0x28ab */
            {8'h00}, /* 0x28aa */
            {8'h00}, /* 0x28a9 */
            {8'h00}, /* 0x28a8 */
            {8'h00}, /* 0x28a7 */
            {8'h00}, /* 0x28a6 */
            {8'h00}, /* 0x28a5 */
            {8'h00}, /* 0x28a4 */
            {8'h00}, /* 0x28a3 */
            {8'h00}, /* 0x28a2 */
            {8'h00}, /* 0x28a1 */
            {8'h00}, /* 0x28a0 */
            {8'h00}, /* 0x289f */
            {8'h00}, /* 0x289e */
            {8'h00}, /* 0x289d */
            {8'h00}, /* 0x289c */
            {8'h00}, /* 0x289b */
            {8'h00}, /* 0x289a */
            {8'h00}, /* 0x2899 */
            {8'h00}, /* 0x2898 */
            {8'h00}, /* 0x2897 */
            {8'h00}, /* 0x2896 */
            {8'h00}, /* 0x2895 */
            {8'h00}, /* 0x2894 */
            {8'h00}, /* 0x2893 */
            {8'h00}, /* 0x2892 */
            {8'h00}, /* 0x2891 */
            {8'h00}, /* 0x2890 */
            {8'h00}, /* 0x288f */
            {8'h00}, /* 0x288e */
            {8'h00}, /* 0x288d */
            {8'h00}, /* 0x288c */
            {8'h00}, /* 0x288b */
            {8'h00}, /* 0x288a */
            {8'h00}, /* 0x2889 */
            {8'h00}, /* 0x2888 */
            {8'h00}, /* 0x2887 */
            {8'h00}, /* 0x2886 */
            {8'h00}, /* 0x2885 */
            {8'h00}, /* 0x2884 */
            {8'h00}, /* 0x2883 */
            {8'h00}, /* 0x2882 */
            {8'h00}, /* 0x2881 */
            {8'h00}, /* 0x2880 */
            {8'h00}, /* 0x287f */
            {8'h00}, /* 0x287e */
            {8'h00}, /* 0x287d */
            {8'h00}, /* 0x287c */
            {8'h00}, /* 0x287b */
            {8'h00}, /* 0x287a */
            {8'h00}, /* 0x2879 */
            {8'h00}, /* 0x2878 */
            {8'h00}, /* 0x2877 */
            {8'h00}, /* 0x2876 */
            {8'h00}, /* 0x2875 */
            {8'h00}, /* 0x2874 */
            {8'h00}, /* 0x2873 */
            {8'h00}, /* 0x2872 */
            {8'h00}, /* 0x2871 */
            {8'h00}, /* 0x2870 */
            {8'h00}, /* 0x286f */
            {8'h00}, /* 0x286e */
            {8'h00}, /* 0x286d */
            {8'h00}, /* 0x286c */
            {8'h00}, /* 0x286b */
            {8'h00}, /* 0x286a */
            {8'h00}, /* 0x2869 */
            {8'h00}, /* 0x2868 */
            {8'h00}, /* 0x2867 */
            {8'h00}, /* 0x2866 */
            {8'h00}, /* 0x2865 */
            {8'h00}, /* 0x2864 */
            {8'h00}, /* 0x2863 */
            {8'h00}, /* 0x2862 */
            {8'h00}, /* 0x2861 */
            {8'h00}, /* 0x2860 */
            {8'h00}, /* 0x285f */
            {8'h00}, /* 0x285e */
            {8'h00}, /* 0x285d */
            {8'h00}, /* 0x285c */
            {8'h00}, /* 0x285b */
            {8'h00}, /* 0x285a */
            {8'h00}, /* 0x2859 */
            {8'h00}, /* 0x2858 */
            {8'h00}, /* 0x2857 */
            {8'h00}, /* 0x2856 */
            {8'h00}, /* 0x2855 */
            {8'h00}, /* 0x2854 */
            {8'h00}, /* 0x2853 */
            {8'h00}, /* 0x2852 */
            {8'h00}, /* 0x2851 */
            {8'h00}, /* 0x2850 */
            {8'h00}, /* 0x284f */
            {8'h00}, /* 0x284e */
            {8'h00}, /* 0x284d */
            {8'h00}, /* 0x284c */
            {8'h00}, /* 0x284b */
            {8'h00}, /* 0x284a */
            {8'h00}, /* 0x2849 */
            {8'h00}, /* 0x2848 */
            {8'h00}, /* 0x2847 */
            {8'h00}, /* 0x2846 */
            {8'h00}, /* 0x2845 */
            {8'h00}, /* 0x2844 */
            {8'h00}, /* 0x2843 */
            {8'h00}, /* 0x2842 */
            {8'h00}, /* 0x2841 */
            {8'h00}, /* 0x2840 */
            {8'h00}, /* 0x283f */
            {8'h00}, /* 0x283e */
            {8'h00}, /* 0x283d */
            {8'h00}, /* 0x283c */
            {8'h00}, /* 0x283b */
            {8'h00}, /* 0x283a */
            {8'h00}, /* 0x2839 */
            {8'h00}, /* 0x2838 */
            {8'h00}, /* 0x2837 */
            {8'h00}, /* 0x2836 */
            {8'h00}, /* 0x2835 */
            {8'h00}, /* 0x2834 */
            {8'h00}, /* 0x2833 */
            {8'h00}, /* 0x2832 */
            {8'h00}, /* 0x2831 */
            {8'h00}, /* 0x2830 */
            {8'h00}, /* 0x282f */
            {8'h00}, /* 0x282e */
            {8'h00}, /* 0x282d */
            {8'h00}, /* 0x282c */
            {8'h00}, /* 0x282b */
            {8'h00}, /* 0x282a */
            {8'h00}, /* 0x2829 */
            {8'h00}, /* 0x2828 */
            {8'h00}, /* 0x2827 */
            {8'h00}, /* 0x2826 */
            {8'h00}, /* 0x2825 */
            {8'h00}, /* 0x2824 */
            {8'h00}, /* 0x2823 */
            {8'h00}, /* 0x2822 */
            {8'h00}, /* 0x2821 */
            {8'h00}, /* 0x2820 */
            {8'h00}, /* 0x281f */
            {8'h00}, /* 0x281e */
            {8'h00}, /* 0x281d */
            {8'h00}, /* 0x281c */
            {8'h00}, /* 0x281b */
            {8'h00}, /* 0x281a */
            {8'h00}, /* 0x2819 */
            {8'h00}, /* 0x2818 */
            {8'h00}, /* 0x2817 */
            {8'h00}, /* 0x2816 */
            {8'h00}, /* 0x2815 */
            {8'h00}, /* 0x2814 */
            {8'h00}, /* 0x2813 */
            {8'h00}, /* 0x2812 */
            {8'h00}, /* 0x2811 */
            {8'h00}, /* 0x2810 */
            {8'h00}, /* 0x280f */
            {8'h00}, /* 0x280e */
            {8'h00}, /* 0x280d */
            {8'h00}, /* 0x280c */
            {8'h00}, /* 0x280b */
            {8'h00}, /* 0x280a */
            {8'h00}, /* 0x2809 */
            {8'h00}, /* 0x2808 */
            {8'h00}, /* 0x2807 */
            {8'h00}, /* 0x2806 */
            {8'h00}, /* 0x2805 */
            {8'h00}, /* 0x2804 */
            {8'h00}, /* 0x2803 */
            {8'h00}, /* 0x2802 */
            {8'h00}, /* 0x2801 */
            {8'h00}, /* 0x2800 */
            {8'h00}, /* 0x27ff */
            {8'h00}, /* 0x27fe */
            {8'h00}, /* 0x27fd */
            {8'h00}, /* 0x27fc */
            {8'h00}, /* 0x27fb */
            {8'h00}, /* 0x27fa */
            {8'h00}, /* 0x27f9 */
            {8'h00}, /* 0x27f8 */
            {8'h00}, /* 0x27f7 */
            {8'h00}, /* 0x27f6 */
            {8'h00}, /* 0x27f5 */
            {8'h00}, /* 0x27f4 */
            {8'h00}, /* 0x27f3 */
            {8'h00}, /* 0x27f2 */
            {8'h00}, /* 0x27f1 */
            {8'h00}, /* 0x27f0 */
            {8'h00}, /* 0x27ef */
            {8'h00}, /* 0x27ee */
            {8'h00}, /* 0x27ed */
            {8'h00}, /* 0x27ec */
            {8'h00}, /* 0x27eb */
            {8'h00}, /* 0x27ea */
            {8'h00}, /* 0x27e9 */
            {8'h00}, /* 0x27e8 */
            {8'h00}, /* 0x27e7 */
            {8'h00}, /* 0x27e6 */
            {8'h00}, /* 0x27e5 */
            {8'h00}, /* 0x27e4 */
            {8'h00}, /* 0x27e3 */
            {8'h00}, /* 0x27e2 */
            {8'h00}, /* 0x27e1 */
            {8'h00}, /* 0x27e0 */
            {8'h00}, /* 0x27df */
            {8'h00}, /* 0x27de */
            {8'h00}, /* 0x27dd */
            {8'h00}, /* 0x27dc */
            {8'h00}, /* 0x27db */
            {8'h00}, /* 0x27da */
            {8'h00}, /* 0x27d9 */
            {8'h00}, /* 0x27d8 */
            {8'h00}, /* 0x27d7 */
            {8'h00}, /* 0x27d6 */
            {8'h00}, /* 0x27d5 */
            {8'h00}, /* 0x27d4 */
            {8'h00}, /* 0x27d3 */
            {8'h00}, /* 0x27d2 */
            {8'h00}, /* 0x27d1 */
            {8'h00}, /* 0x27d0 */
            {8'h00}, /* 0x27cf */
            {8'h00}, /* 0x27ce */
            {8'h00}, /* 0x27cd */
            {8'h00}, /* 0x27cc */
            {8'h00}, /* 0x27cb */
            {8'h00}, /* 0x27ca */
            {8'h00}, /* 0x27c9 */
            {8'h00}, /* 0x27c8 */
            {8'h00}, /* 0x27c7 */
            {8'h00}, /* 0x27c6 */
            {8'h00}, /* 0x27c5 */
            {8'h00}, /* 0x27c4 */
            {8'h00}, /* 0x27c3 */
            {8'h00}, /* 0x27c2 */
            {8'h00}, /* 0x27c1 */
            {8'h00}, /* 0x27c0 */
            {8'h00}, /* 0x27bf */
            {8'h00}, /* 0x27be */
            {8'h00}, /* 0x27bd */
            {8'h00}, /* 0x27bc */
            {8'h00}, /* 0x27bb */
            {8'h00}, /* 0x27ba */
            {8'h00}, /* 0x27b9 */
            {8'h00}, /* 0x27b8 */
            {8'h00}, /* 0x27b7 */
            {8'h00}, /* 0x27b6 */
            {8'h00}, /* 0x27b5 */
            {8'h00}, /* 0x27b4 */
            {8'h00}, /* 0x27b3 */
            {8'h00}, /* 0x27b2 */
            {8'h00}, /* 0x27b1 */
            {8'h00}, /* 0x27b0 */
            {8'h00}, /* 0x27af */
            {8'h00}, /* 0x27ae */
            {8'h00}, /* 0x27ad */
            {8'h00}, /* 0x27ac */
            {8'h00}, /* 0x27ab */
            {8'h00}, /* 0x27aa */
            {8'h00}, /* 0x27a9 */
            {8'h00}, /* 0x27a8 */
            {8'h00}, /* 0x27a7 */
            {8'h00}, /* 0x27a6 */
            {8'h00}, /* 0x27a5 */
            {8'h00}, /* 0x27a4 */
            {8'h00}, /* 0x27a3 */
            {8'h00}, /* 0x27a2 */
            {8'h00}, /* 0x27a1 */
            {8'h00}, /* 0x27a0 */
            {8'h00}, /* 0x279f */
            {8'h00}, /* 0x279e */
            {8'h00}, /* 0x279d */
            {8'h00}, /* 0x279c */
            {8'h00}, /* 0x279b */
            {8'h00}, /* 0x279a */
            {8'h00}, /* 0x2799 */
            {8'h00}, /* 0x2798 */
            {8'h00}, /* 0x2797 */
            {8'h00}, /* 0x2796 */
            {8'h00}, /* 0x2795 */
            {8'h00}, /* 0x2794 */
            {8'h00}, /* 0x2793 */
            {8'h00}, /* 0x2792 */
            {8'h00}, /* 0x2791 */
            {8'h00}, /* 0x2790 */
            {8'h00}, /* 0x278f */
            {8'h00}, /* 0x278e */
            {8'h00}, /* 0x278d */
            {8'h00}, /* 0x278c */
            {8'h00}, /* 0x278b */
            {8'h00}, /* 0x278a */
            {8'h00}, /* 0x2789 */
            {8'h00}, /* 0x2788 */
            {8'h00}, /* 0x2787 */
            {8'h00}, /* 0x2786 */
            {8'h00}, /* 0x2785 */
            {8'h00}, /* 0x2784 */
            {8'h00}, /* 0x2783 */
            {8'h00}, /* 0x2782 */
            {8'h00}, /* 0x2781 */
            {8'h00}, /* 0x2780 */
            {8'h00}, /* 0x277f */
            {8'h00}, /* 0x277e */
            {8'h00}, /* 0x277d */
            {8'h00}, /* 0x277c */
            {8'h00}, /* 0x277b */
            {8'h00}, /* 0x277a */
            {8'h00}, /* 0x2779 */
            {8'h00}, /* 0x2778 */
            {8'h00}, /* 0x2777 */
            {8'h00}, /* 0x2776 */
            {8'h00}, /* 0x2775 */
            {8'h00}, /* 0x2774 */
            {8'h00}, /* 0x2773 */
            {8'h00}, /* 0x2772 */
            {8'h00}, /* 0x2771 */
            {8'h00}, /* 0x2770 */
            {8'h00}, /* 0x276f */
            {8'h00}, /* 0x276e */
            {8'h00}, /* 0x276d */
            {8'h00}, /* 0x276c */
            {8'h00}, /* 0x276b */
            {8'h00}, /* 0x276a */
            {8'h00}, /* 0x2769 */
            {8'h00}, /* 0x2768 */
            {8'h00}, /* 0x2767 */
            {8'h00}, /* 0x2766 */
            {8'h00}, /* 0x2765 */
            {8'h00}, /* 0x2764 */
            {8'h00}, /* 0x2763 */
            {8'h00}, /* 0x2762 */
            {8'h00}, /* 0x2761 */
            {8'h00}, /* 0x2760 */
            {8'h00}, /* 0x275f */
            {8'h00}, /* 0x275e */
            {8'h00}, /* 0x275d */
            {8'h00}, /* 0x275c */
            {8'h00}, /* 0x275b */
            {8'h00}, /* 0x275a */
            {8'h00}, /* 0x2759 */
            {8'h00}, /* 0x2758 */
            {8'h00}, /* 0x2757 */
            {8'h00}, /* 0x2756 */
            {8'h00}, /* 0x2755 */
            {8'h00}, /* 0x2754 */
            {8'h00}, /* 0x2753 */
            {8'h00}, /* 0x2752 */
            {8'h00}, /* 0x2751 */
            {8'h00}, /* 0x2750 */
            {8'h00}, /* 0x274f */
            {8'h00}, /* 0x274e */
            {8'h00}, /* 0x274d */
            {8'h00}, /* 0x274c */
            {8'h00}, /* 0x274b */
            {8'h00}, /* 0x274a */
            {8'h00}, /* 0x2749 */
            {8'h00}, /* 0x2748 */
            {8'h00}, /* 0x2747 */
            {8'h00}, /* 0x2746 */
            {8'h00}, /* 0x2745 */
            {8'h00}, /* 0x2744 */
            {8'h00}, /* 0x2743 */
            {8'h00}, /* 0x2742 */
            {8'h00}, /* 0x2741 */
            {8'h00}, /* 0x2740 */
            {8'h00}, /* 0x273f */
            {8'h00}, /* 0x273e */
            {8'h00}, /* 0x273d */
            {8'h00}, /* 0x273c */
            {8'h00}, /* 0x273b */
            {8'h00}, /* 0x273a */
            {8'h00}, /* 0x2739 */
            {8'h00}, /* 0x2738 */
            {8'h00}, /* 0x2737 */
            {8'h00}, /* 0x2736 */
            {8'h00}, /* 0x2735 */
            {8'h00}, /* 0x2734 */
            {8'h00}, /* 0x2733 */
            {8'h00}, /* 0x2732 */
            {8'h00}, /* 0x2731 */
            {8'h00}, /* 0x2730 */
            {8'h00}, /* 0x272f */
            {8'h00}, /* 0x272e */
            {8'h00}, /* 0x272d */
            {8'h00}, /* 0x272c */
            {8'h00}, /* 0x272b */
            {8'h00}, /* 0x272a */
            {8'h00}, /* 0x2729 */
            {8'h00}, /* 0x2728 */
            {8'h00}, /* 0x2727 */
            {8'h00}, /* 0x2726 */
            {8'h00}, /* 0x2725 */
            {8'h00}, /* 0x2724 */
            {8'h00}, /* 0x2723 */
            {8'h00}, /* 0x2722 */
            {8'h00}, /* 0x2721 */
            {8'h00}, /* 0x2720 */
            {8'h00}, /* 0x271f */
            {8'h00}, /* 0x271e */
            {8'h00}, /* 0x271d */
            {8'h00}, /* 0x271c */
            {8'h00}, /* 0x271b */
            {8'h00}, /* 0x271a */
            {8'h00}, /* 0x2719 */
            {8'h00}, /* 0x2718 */
            {8'h00}, /* 0x2717 */
            {8'h00}, /* 0x2716 */
            {8'h00}, /* 0x2715 */
            {8'h00}, /* 0x2714 */
            {8'h00}, /* 0x2713 */
            {8'h00}, /* 0x2712 */
            {8'h00}, /* 0x2711 */
            {8'h00}, /* 0x2710 */
            {8'h00}, /* 0x270f */
            {8'h00}, /* 0x270e */
            {8'h00}, /* 0x270d */
            {8'h00}, /* 0x270c */
            {8'h00}, /* 0x270b */
            {8'h00}, /* 0x270a */
            {8'h00}, /* 0x2709 */
            {8'h00}, /* 0x2708 */
            {8'h00}, /* 0x2707 */
            {8'h00}, /* 0x2706 */
            {8'h00}, /* 0x2705 */
            {8'h00}, /* 0x2704 */
            {8'h00}, /* 0x2703 */
            {8'h00}, /* 0x2702 */
            {8'h00}, /* 0x2701 */
            {8'h00}, /* 0x2700 */
            {8'h00}, /* 0x26ff */
            {8'h00}, /* 0x26fe */
            {8'h00}, /* 0x26fd */
            {8'h00}, /* 0x26fc */
            {8'h00}, /* 0x26fb */
            {8'h00}, /* 0x26fa */
            {8'h00}, /* 0x26f9 */
            {8'h00}, /* 0x26f8 */
            {8'h00}, /* 0x26f7 */
            {8'h00}, /* 0x26f6 */
            {8'h00}, /* 0x26f5 */
            {8'h00}, /* 0x26f4 */
            {8'h00}, /* 0x26f3 */
            {8'h00}, /* 0x26f2 */
            {8'h00}, /* 0x26f1 */
            {8'h00}, /* 0x26f0 */
            {8'h00}, /* 0x26ef */
            {8'h00}, /* 0x26ee */
            {8'h00}, /* 0x26ed */
            {8'h00}, /* 0x26ec */
            {8'h00}, /* 0x26eb */
            {8'h00}, /* 0x26ea */
            {8'h00}, /* 0x26e9 */
            {8'h00}, /* 0x26e8 */
            {8'h00}, /* 0x26e7 */
            {8'h00}, /* 0x26e6 */
            {8'h00}, /* 0x26e5 */
            {8'h00}, /* 0x26e4 */
            {8'h00}, /* 0x26e3 */
            {8'h00}, /* 0x26e2 */
            {8'h00}, /* 0x26e1 */
            {8'h00}, /* 0x26e0 */
            {8'h00}, /* 0x26df */
            {8'h00}, /* 0x26de */
            {8'h00}, /* 0x26dd */
            {8'h00}, /* 0x26dc */
            {8'h00}, /* 0x26db */
            {8'h00}, /* 0x26da */
            {8'h00}, /* 0x26d9 */
            {8'h00}, /* 0x26d8 */
            {8'h00}, /* 0x26d7 */
            {8'h00}, /* 0x26d6 */
            {8'h00}, /* 0x26d5 */
            {8'h00}, /* 0x26d4 */
            {8'h00}, /* 0x26d3 */
            {8'h00}, /* 0x26d2 */
            {8'h00}, /* 0x26d1 */
            {8'h00}, /* 0x26d0 */
            {8'h00}, /* 0x26cf */
            {8'h00}, /* 0x26ce */
            {8'h00}, /* 0x26cd */
            {8'h00}, /* 0x26cc */
            {8'h00}, /* 0x26cb */
            {8'h00}, /* 0x26ca */
            {8'h00}, /* 0x26c9 */
            {8'h00}, /* 0x26c8 */
            {8'h00}, /* 0x26c7 */
            {8'h00}, /* 0x26c6 */
            {8'h00}, /* 0x26c5 */
            {8'h00}, /* 0x26c4 */
            {8'h00}, /* 0x26c3 */
            {8'h00}, /* 0x26c2 */
            {8'h00}, /* 0x26c1 */
            {8'h00}, /* 0x26c0 */
            {8'h00}, /* 0x26bf */
            {8'h00}, /* 0x26be */
            {8'h00}, /* 0x26bd */
            {8'h00}, /* 0x26bc */
            {8'h00}, /* 0x26bb */
            {8'h00}, /* 0x26ba */
            {8'h00}, /* 0x26b9 */
            {8'h00}, /* 0x26b8 */
            {8'h00}, /* 0x26b7 */
            {8'h00}, /* 0x26b6 */
            {8'h00}, /* 0x26b5 */
            {8'h00}, /* 0x26b4 */
            {8'h00}, /* 0x26b3 */
            {8'h00}, /* 0x26b2 */
            {8'h00}, /* 0x26b1 */
            {8'h00}, /* 0x26b0 */
            {8'h00}, /* 0x26af */
            {8'h00}, /* 0x26ae */
            {8'h00}, /* 0x26ad */
            {8'h00}, /* 0x26ac */
            {8'h00}, /* 0x26ab */
            {8'h00}, /* 0x26aa */
            {8'h00}, /* 0x26a9 */
            {8'h00}, /* 0x26a8 */
            {8'h00}, /* 0x26a7 */
            {8'h00}, /* 0x26a6 */
            {8'h00}, /* 0x26a5 */
            {8'h00}, /* 0x26a4 */
            {8'h00}, /* 0x26a3 */
            {8'h00}, /* 0x26a2 */
            {8'h00}, /* 0x26a1 */
            {8'h00}, /* 0x26a0 */
            {8'h00}, /* 0x269f */
            {8'h00}, /* 0x269e */
            {8'h00}, /* 0x269d */
            {8'h00}, /* 0x269c */
            {8'h00}, /* 0x269b */
            {8'h00}, /* 0x269a */
            {8'h00}, /* 0x2699 */
            {8'h00}, /* 0x2698 */
            {8'h00}, /* 0x2697 */
            {8'h00}, /* 0x2696 */
            {8'h00}, /* 0x2695 */
            {8'h00}, /* 0x2694 */
            {8'h00}, /* 0x2693 */
            {8'h00}, /* 0x2692 */
            {8'h00}, /* 0x2691 */
            {8'h00}, /* 0x2690 */
            {8'h00}, /* 0x268f */
            {8'h00}, /* 0x268e */
            {8'h00}, /* 0x268d */
            {8'h00}, /* 0x268c */
            {8'h00}, /* 0x268b */
            {8'h00}, /* 0x268a */
            {8'h00}, /* 0x2689 */
            {8'h00}, /* 0x2688 */
            {8'h00}, /* 0x2687 */
            {8'h00}, /* 0x2686 */
            {8'h00}, /* 0x2685 */
            {8'h00}, /* 0x2684 */
            {8'h00}, /* 0x2683 */
            {8'h00}, /* 0x2682 */
            {8'h00}, /* 0x2681 */
            {8'h00}, /* 0x2680 */
            {8'h00}, /* 0x267f */
            {8'h00}, /* 0x267e */
            {8'h00}, /* 0x267d */
            {8'h00}, /* 0x267c */
            {8'h00}, /* 0x267b */
            {8'h00}, /* 0x267a */
            {8'h00}, /* 0x2679 */
            {8'h00}, /* 0x2678 */
            {8'h00}, /* 0x2677 */
            {8'h00}, /* 0x2676 */
            {8'h00}, /* 0x2675 */
            {8'h00}, /* 0x2674 */
            {8'h00}, /* 0x2673 */
            {8'h00}, /* 0x2672 */
            {8'h00}, /* 0x2671 */
            {8'h00}, /* 0x2670 */
            {8'h00}, /* 0x266f */
            {8'h00}, /* 0x266e */
            {8'h00}, /* 0x266d */
            {8'h00}, /* 0x266c */
            {8'h00}, /* 0x266b */
            {8'h00}, /* 0x266a */
            {8'h00}, /* 0x2669 */
            {8'h00}, /* 0x2668 */
            {8'h00}, /* 0x2667 */
            {8'h00}, /* 0x2666 */
            {8'h00}, /* 0x2665 */
            {8'h00}, /* 0x2664 */
            {8'h00}, /* 0x2663 */
            {8'h00}, /* 0x2662 */
            {8'h00}, /* 0x2661 */
            {8'h00}, /* 0x2660 */
            {8'h00}, /* 0x265f */
            {8'h00}, /* 0x265e */
            {8'h00}, /* 0x265d */
            {8'h00}, /* 0x265c */
            {8'h00}, /* 0x265b */
            {8'h00}, /* 0x265a */
            {8'h00}, /* 0x2659 */
            {8'h00}, /* 0x2658 */
            {8'h00}, /* 0x2657 */
            {8'h00}, /* 0x2656 */
            {8'h00}, /* 0x2655 */
            {8'h00}, /* 0x2654 */
            {8'h00}, /* 0x2653 */
            {8'h00}, /* 0x2652 */
            {8'h00}, /* 0x2651 */
            {8'h00}, /* 0x2650 */
            {8'h00}, /* 0x264f */
            {8'h00}, /* 0x264e */
            {8'h00}, /* 0x264d */
            {8'h00}, /* 0x264c */
            {8'h00}, /* 0x264b */
            {8'h00}, /* 0x264a */
            {8'h00}, /* 0x2649 */
            {8'h00}, /* 0x2648 */
            {8'h00}, /* 0x2647 */
            {8'h00}, /* 0x2646 */
            {8'h00}, /* 0x2645 */
            {8'h00}, /* 0x2644 */
            {8'h00}, /* 0x2643 */
            {8'h00}, /* 0x2642 */
            {8'h00}, /* 0x2641 */
            {8'h00}, /* 0x2640 */
            {8'h00}, /* 0x263f */
            {8'h00}, /* 0x263e */
            {8'h00}, /* 0x263d */
            {8'h00}, /* 0x263c */
            {8'h00}, /* 0x263b */
            {8'h00}, /* 0x263a */
            {8'h00}, /* 0x2639 */
            {8'h00}, /* 0x2638 */
            {8'h00}, /* 0x2637 */
            {8'h00}, /* 0x2636 */
            {8'h00}, /* 0x2635 */
            {8'h00}, /* 0x2634 */
            {8'h00}, /* 0x2633 */
            {8'h00}, /* 0x2632 */
            {8'h00}, /* 0x2631 */
            {8'h00}, /* 0x2630 */
            {8'h00}, /* 0x262f */
            {8'h00}, /* 0x262e */
            {8'h00}, /* 0x262d */
            {8'h00}, /* 0x262c */
            {8'h00}, /* 0x262b */
            {8'h00}, /* 0x262a */
            {8'h00}, /* 0x2629 */
            {8'h00}, /* 0x2628 */
            {8'h00}, /* 0x2627 */
            {8'h00}, /* 0x2626 */
            {8'h00}, /* 0x2625 */
            {8'h00}, /* 0x2624 */
            {8'h00}, /* 0x2623 */
            {8'h00}, /* 0x2622 */
            {8'h00}, /* 0x2621 */
            {8'h00}, /* 0x2620 */
            {8'h00}, /* 0x261f */
            {8'h00}, /* 0x261e */
            {8'h00}, /* 0x261d */
            {8'h00}, /* 0x261c */
            {8'h00}, /* 0x261b */
            {8'h00}, /* 0x261a */
            {8'h00}, /* 0x2619 */
            {8'h00}, /* 0x2618 */
            {8'h00}, /* 0x2617 */
            {8'h00}, /* 0x2616 */
            {8'h00}, /* 0x2615 */
            {8'h00}, /* 0x2614 */
            {8'h00}, /* 0x2613 */
            {8'h00}, /* 0x2612 */
            {8'h00}, /* 0x2611 */
            {8'h00}, /* 0x2610 */
            {8'h00}, /* 0x260f */
            {8'h00}, /* 0x260e */
            {8'h00}, /* 0x260d */
            {8'h00}, /* 0x260c */
            {8'h00}, /* 0x260b */
            {8'h00}, /* 0x260a */
            {8'h00}, /* 0x2609 */
            {8'h00}, /* 0x2608 */
            {8'h00}, /* 0x2607 */
            {8'h00}, /* 0x2606 */
            {8'h00}, /* 0x2605 */
            {8'h00}, /* 0x2604 */
            {8'h00}, /* 0x2603 */
            {8'h00}, /* 0x2602 */
            {8'h00}, /* 0x2601 */
            {8'h00}, /* 0x2600 */
            {8'h00}, /* 0x25ff */
            {8'h00}, /* 0x25fe */
            {8'h00}, /* 0x25fd */
            {8'h00}, /* 0x25fc */
            {8'h00}, /* 0x25fb */
            {8'h00}, /* 0x25fa */
            {8'h00}, /* 0x25f9 */
            {8'h00}, /* 0x25f8 */
            {8'h00}, /* 0x25f7 */
            {8'h00}, /* 0x25f6 */
            {8'h00}, /* 0x25f5 */
            {8'h00}, /* 0x25f4 */
            {8'h00}, /* 0x25f3 */
            {8'h00}, /* 0x25f2 */
            {8'h00}, /* 0x25f1 */
            {8'h00}, /* 0x25f0 */
            {8'h00}, /* 0x25ef */
            {8'h00}, /* 0x25ee */
            {8'h00}, /* 0x25ed */
            {8'h00}, /* 0x25ec */
            {8'h00}, /* 0x25eb */
            {8'h00}, /* 0x25ea */
            {8'h00}, /* 0x25e9 */
            {8'h00}, /* 0x25e8 */
            {8'h00}, /* 0x25e7 */
            {8'h00}, /* 0x25e6 */
            {8'h00}, /* 0x25e5 */
            {8'h00}, /* 0x25e4 */
            {8'h00}, /* 0x25e3 */
            {8'h00}, /* 0x25e2 */
            {8'h00}, /* 0x25e1 */
            {8'h00}, /* 0x25e0 */
            {8'h00}, /* 0x25df */
            {8'h00}, /* 0x25de */
            {8'h00}, /* 0x25dd */
            {8'h00}, /* 0x25dc */
            {8'h00}, /* 0x25db */
            {8'h00}, /* 0x25da */
            {8'h00}, /* 0x25d9 */
            {8'h00}, /* 0x25d8 */
            {8'h00}, /* 0x25d7 */
            {8'h00}, /* 0x25d6 */
            {8'h00}, /* 0x25d5 */
            {8'h00}, /* 0x25d4 */
            {8'h00}, /* 0x25d3 */
            {8'h00}, /* 0x25d2 */
            {8'h00}, /* 0x25d1 */
            {8'h00}, /* 0x25d0 */
            {8'h00}, /* 0x25cf */
            {8'h00}, /* 0x25ce */
            {8'h00}, /* 0x25cd */
            {8'h00}, /* 0x25cc */
            {8'h00}, /* 0x25cb */
            {8'h00}, /* 0x25ca */
            {8'h00}, /* 0x25c9 */
            {8'h00}, /* 0x25c8 */
            {8'h00}, /* 0x25c7 */
            {8'h00}, /* 0x25c6 */
            {8'h00}, /* 0x25c5 */
            {8'h00}, /* 0x25c4 */
            {8'h00}, /* 0x25c3 */
            {8'h00}, /* 0x25c2 */
            {8'h00}, /* 0x25c1 */
            {8'h00}, /* 0x25c0 */
            {8'h00}, /* 0x25bf */
            {8'h00}, /* 0x25be */
            {8'h00}, /* 0x25bd */
            {8'h00}, /* 0x25bc */
            {8'h00}, /* 0x25bb */
            {8'h00}, /* 0x25ba */
            {8'h00}, /* 0x25b9 */
            {8'h00}, /* 0x25b8 */
            {8'h00}, /* 0x25b7 */
            {8'h00}, /* 0x25b6 */
            {8'h00}, /* 0x25b5 */
            {8'h00}, /* 0x25b4 */
            {8'h00}, /* 0x25b3 */
            {8'h00}, /* 0x25b2 */
            {8'h00}, /* 0x25b1 */
            {8'h00}, /* 0x25b0 */
            {8'h00}, /* 0x25af */
            {8'h00}, /* 0x25ae */
            {8'h00}, /* 0x25ad */
            {8'h00}, /* 0x25ac */
            {8'h00}, /* 0x25ab */
            {8'h00}, /* 0x25aa */
            {8'h00}, /* 0x25a9 */
            {8'h00}, /* 0x25a8 */
            {8'h00}, /* 0x25a7 */
            {8'h00}, /* 0x25a6 */
            {8'h00}, /* 0x25a5 */
            {8'h00}, /* 0x25a4 */
            {8'h00}, /* 0x25a3 */
            {8'h00}, /* 0x25a2 */
            {8'h00}, /* 0x25a1 */
            {8'h00}, /* 0x25a0 */
            {8'h00}, /* 0x259f */
            {8'h00}, /* 0x259e */
            {8'h00}, /* 0x259d */
            {8'h00}, /* 0x259c */
            {8'h00}, /* 0x259b */
            {8'h00}, /* 0x259a */
            {8'h00}, /* 0x2599 */
            {8'h00}, /* 0x2598 */
            {8'h00}, /* 0x2597 */
            {8'h00}, /* 0x2596 */
            {8'h00}, /* 0x2595 */
            {8'h00}, /* 0x2594 */
            {8'h00}, /* 0x2593 */
            {8'h00}, /* 0x2592 */
            {8'h00}, /* 0x2591 */
            {8'h00}, /* 0x2590 */
            {8'h00}, /* 0x258f */
            {8'h00}, /* 0x258e */
            {8'h00}, /* 0x258d */
            {8'h00}, /* 0x258c */
            {8'h00}, /* 0x258b */
            {8'h00}, /* 0x258a */
            {8'h00}, /* 0x2589 */
            {8'h00}, /* 0x2588 */
            {8'h00}, /* 0x2587 */
            {8'h00}, /* 0x2586 */
            {8'h00}, /* 0x2585 */
            {8'h00}, /* 0x2584 */
            {8'h00}, /* 0x2583 */
            {8'h00}, /* 0x2582 */
            {8'h00}, /* 0x2581 */
            {8'h00}, /* 0x2580 */
            {8'h00}, /* 0x257f */
            {8'h00}, /* 0x257e */
            {8'h00}, /* 0x257d */
            {8'h00}, /* 0x257c */
            {8'h00}, /* 0x257b */
            {8'h00}, /* 0x257a */
            {8'h00}, /* 0x2579 */
            {8'h00}, /* 0x2578 */
            {8'h00}, /* 0x2577 */
            {8'h00}, /* 0x2576 */
            {8'h00}, /* 0x2575 */
            {8'h00}, /* 0x2574 */
            {8'h00}, /* 0x2573 */
            {8'h00}, /* 0x2572 */
            {8'h00}, /* 0x2571 */
            {8'h00}, /* 0x2570 */
            {8'h00}, /* 0x256f */
            {8'h00}, /* 0x256e */
            {8'h00}, /* 0x256d */
            {8'h00}, /* 0x256c */
            {8'h00}, /* 0x256b */
            {8'h00}, /* 0x256a */
            {8'h00}, /* 0x2569 */
            {8'h00}, /* 0x2568 */
            {8'h00}, /* 0x2567 */
            {8'h00}, /* 0x2566 */
            {8'h00}, /* 0x2565 */
            {8'h00}, /* 0x2564 */
            {8'h00}, /* 0x2563 */
            {8'h00}, /* 0x2562 */
            {8'h00}, /* 0x2561 */
            {8'h00}, /* 0x2560 */
            {8'h00}, /* 0x255f */
            {8'h00}, /* 0x255e */
            {8'h00}, /* 0x255d */
            {8'h00}, /* 0x255c */
            {8'h00}, /* 0x255b */
            {8'h00}, /* 0x255a */
            {8'h00}, /* 0x2559 */
            {8'h00}, /* 0x2558 */
            {8'h00}, /* 0x2557 */
            {8'h00}, /* 0x2556 */
            {8'h00}, /* 0x2555 */
            {8'h00}, /* 0x2554 */
            {8'h00}, /* 0x2553 */
            {8'h00}, /* 0x2552 */
            {8'h00}, /* 0x2551 */
            {8'h00}, /* 0x2550 */
            {8'h00}, /* 0x254f */
            {8'h00}, /* 0x254e */
            {8'h00}, /* 0x254d */
            {8'h00}, /* 0x254c */
            {8'h00}, /* 0x254b */
            {8'h00}, /* 0x254a */
            {8'h00}, /* 0x2549 */
            {8'h00}, /* 0x2548 */
            {8'h00}, /* 0x2547 */
            {8'h00}, /* 0x2546 */
            {8'h00}, /* 0x2545 */
            {8'h00}, /* 0x2544 */
            {8'h00}, /* 0x2543 */
            {8'h00}, /* 0x2542 */
            {8'h00}, /* 0x2541 */
            {8'h00}, /* 0x2540 */
            {8'h00}, /* 0x253f */
            {8'h00}, /* 0x253e */
            {8'h00}, /* 0x253d */
            {8'h00}, /* 0x253c */
            {8'h00}, /* 0x253b */
            {8'h00}, /* 0x253a */
            {8'h00}, /* 0x2539 */
            {8'h00}, /* 0x2538 */
            {8'h00}, /* 0x2537 */
            {8'h00}, /* 0x2536 */
            {8'h00}, /* 0x2535 */
            {8'h00}, /* 0x2534 */
            {8'h00}, /* 0x2533 */
            {8'h00}, /* 0x2532 */
            {8'h00}, /* 0x2531 */
            {8'h00}, /* 0x2530 */
            {8'h00}, /* 0x252f */
            {8'h00}, /* 0x252e */
            {8'h00}, /* 0x252d */
            {8'h00}, /* 0x252c */
            {8'h00}, /* 0x252b */
            {8'h00}, /* 0x252a */
            {8'h00}, /* 0x2529 */
            {8'h00}, /* 0x2528 */
            {8'h00}, /* 0x2527 */
            {8'h00}, /* 0x2526 */
            {8'h00}, /* 0x2525 */
            {8'h00}, /* 0x2524 */
            {8'h00}, /* 0x2523 */
            {8'h00}, /* 0x2522 */
            {8'h00}, /* 0x2521 */
            {8'h00}, /* 0x2520 */
            {8'h00}, /* 0x251f */
            {8'h00}, /* 0x251e */
            {8'h00}, /* 0x251d */
            {8'h00}, /* 0x251c */
            {8'h00}, /* 0x251b */
            {8'h00}, /* 0x251a */
            {8'h00}, /* 0x2519 */
            {8'h00}, /* 0x2518 */
            {8'h00}, /* 0x2517 */
            {8'h00}, /* 0x2516 */
            {8'h00}, /* 0x2515 */
            {8'h00}, /* 0x2514 */
            {8'h00}, /* 0x2513 */
            {8'h00}, /* 0x2512 */
            {8'h00}, /* 0x2511 */
            {8'h00}, /* 0x2510 */
            {8'h00}, /* 0x250f */
            {8'h00}, /* 0x250e */
            {8'h00}, /* 0x250d */
            {8'h00}, /* 0x250c */
            {8'h00}, /* 0x250b */
            {8'h00}, /* 0x250a */
            {8'h00}, /* 0x2509 */
            {8'h00}, /* 0x2508 */
            {8'h00}, /* 0x2507 */
            {8'h00}, /* 0x2506 */
            {8'h00}, /* 0x2505 */
            {8'h00}, /* 0x2504 */
            {8'h00}, /* 0x2503 */
            {8'h00}, /* 0x2502 */
            {8'h00}, /* 0x2501 */
            {8'h00}, /* 0x2500 */
            {8'h00}, /* 0x24ff */
            {8'h00}, /* 0x24fe */
            {8'h00}, /* 0x24fd */
            {8'h00}, /* 0x24fc */
            {8'h00}, /* 0x24fb */
            {8'h00}, /* 0x24fa */
            {8'h00}, /* 0x24f9 */
            {8'h00}, /* 0x24f8 */
            {8'h00}, /* 0x24f7 */
            {8'h00}, /* 0x24f6 */
            {8'h00}, /* 0x24f5 */
            {8'h00}, /* 0x24f4 */
            {8'h00}, /* 0x24f3 */
            {8'h00}, /* 0x24f2 */
            {8'h00}, /* 0x24f1 */
            {8'h00}, /* 0x24f0 */
            {8'h00}, /* 0x24ef */
            {8'h00}, /* 0x24ee */
            {8'h00}, /* 0x24ed */
            {8'h00}, /* 0x24ec */
            {8'h00}, /* 0x24eb */
            {8'h00}, /* 0x24ea */
            {8'h00}, /* 0x24e9 */
            {8'h00}, /* 0x24e8 */
            {8'h00}, /* 0x24e7 */
            {8'h00}, /* 0x24e6 */
            {8'h00}, /* 0x24e5 */
            {8'h00}, /* 0x24e4 */
            {8'h00}, /* 0x24e3 */
            {8'h00}, /* 0x24e2 */
            {8'h00}, /* 0x24e1 */
            {8'h00}, /* 0x24e0 */
            {8'h00}, /* 0x24df */
            {8'h00}, /* 0x24de */
            {8'h00}, /* 0x24dd */
            {8'h00}, /* 0x24dc */
            {8'h00}, /* 0x24db */
            {8'h00}, /* 0x24da */
            {8'h00}, /* 0x24d9 */
            {8'h00}, /* 0x24d8 */
            {8'h00}, /* 0x24d7 */
            {8'h00}, /* 0x24d6 */
            {8'h00}, /* 0x24d5 */
            {8'h00}, /* 0x24d4 */
            {8'h00}, /* 0x24d3 */
            {8'h00}, /* 0x24d2 */
            {8'h00}, /* 0x24d1 */
            {8'h00}, /* 0x24d0 */
            {8'h00}, /* 0x24cf */
            {8'h00}, /* 0x24ce */
            {8'h00}, /* 0x24cd */
            {8'h00}, /* 0x24cc */
            {8'h00}, /* 0x24cb */
            {8'h00}, /* 0x24ca */
            {8'h00}, /* 0x24c9 */
            {8'h00}, /* 0x24c8 */
            {8'h00}, /* 0x24c7 */
            {8'h00}, /* 0x24c6 */
            {8'h00}, /* 0x24c5 */
            {8'h00}, /* 0x24c4 */
            {8'h00}, /* 0x24c3 */
            {8'h00}, /* 0x24c2 */
            {8'h00}, /* 0x24c1 */
            {8'h00}, /* 0x24c0 */
            {8'h00}, /* 0x24bf */
            {8'h00}, /* 0x24be */
            {8'h00}, /* 0x24bd */
            {8'h00}, /* 0x24bc */
            {8'h00}, /* 0x24bb */
            {8'h00}, /* 0x24ba */
            {8'h00}, /* 0x24b9 */
            {8'h00}, /* 0x24b8 */
            {8'h00}, /* 0x24b7 */
            {8'h00}, /* 0x24b6 */
            {8'h00}, /* 0x24b5 */
            {8'h00}, /* 0x24b4 */
            {8'h00}, /* 0x24b3 */
            {8'h00}, /* 0x24b2 */
            {8'h00}, /* 0x24b1 */
            {8'h00}, /* 0x24b0 */
            {8'h00}, /* 0x24af */
            {8'h00}, /* 0x24ae */
            {8'h00}, /* 0x24ad */
            {8'h00}, /* 0x24ac */
            {8'h00}, /* 0x24ab */
            {8'h00}, /* 0x24aa */
            {8'h00}, /* 0x24a9 */
            {8'h00}, /* 0x24a8 */
            {8'h00}, /* 0x24a7 */
            {8'h00}, /* 0x24a6 */
            {8'h00}, /* 0x24a5 */
            {8'h00}, /* 0x24a4 */
            {8'h00}, /* 0x24a3 */
            {8'h00}, /* 0x24a2 */
            {8'h00}, /* 0x24a1 */
            {8'h00}, /* 0x24a0 */
            {8'h00}, /* 0x249f */
            {8'h00}, /* 0x249e */
            {8'h00}, /* 0x249d */
            {8'h00}, /* 0x249c */
            {8'h00}, /* 0x249b */
            {8'h00}, /* 0x249a */
            {8'h00}, /* 0x2499 */
            {8'h00}, /* 0x2498 */
            {8'h00}, /* 0x2497 */
            {8'h00}, /* 0x2496 */
            {8'h00}, /* 0x2495 */
            {8'h00}, /* 0x2494 */
            {8'h00}, /* 0x2493 */
            {8'h00}, /* 0x2492 */
            {8'h00}, /* 0x2491 */
            {8'h00}, /* 0x2490 */
            {8'h00}, /* 0x248f */
            {8'h00}, /* 0x248e */
            {8'h00}, /* 0x248d */
            {8'h00}, /* 0x248c */
            {8'h00}, /* 0x248b */
            {8'h00}, /* 0x248a */
            {8'h00}, /* 0x2489 */
            {8'h00}, /* 0x2488 */
            {8'h00}, /* 0x2487 */
            {8'h00}, /* 0x2486 */
            {8'h00}, /* 0x2485 */
            {8'h00}, /* 0x2484 */
            {8'h00}, /* 0x2483 */
            {8'h00}, /* 0x2482 */
            {8'h00}, /* 0x2481 */
            {8'h00}, /* 0x2480 */
            {8'h00}, /* 0x247f */
            {8'h00}, /* 0x247e */
            {8'h00}, /* 0x247d */
            {8'h00}, /* 0x247c */
            {8'h00}, /* 0x247b */
            {8'h00}, /* 0x247a */
            {8'h00}, /* 0x2479 */
            {8'h00}, /* 0x2478 */
            {8'h00}, /* 0x2477 */
            {8'h00}, /* 0x2476 */
            {8'h00}, /* 0x2475 */
            {8'h00}, /* 0x2474 */
            {8'h00}, /* 0x2473 */
            {8'h00}, /* 0x2472 */
            {8'h00}, /* 0x2471 */
            {8'h00}, /* 0x2470 */
            {8'h00}, /* 0x246f */
            {8'h00}, /* 0x246e */
            {8'h00}, /* 0x246d */
            {8'h00}, /* 0x246c */
            {8'h00}, /* 0x246b */
            {8'h00}, /* 0x246a */
            {8'h00}, /* 0x2469 */
            {8'h00}, /* 0x2468 */
            {8'h00}, /* 0x2467 */
            {8'h00}, /* 0x2466 */
            {8'h00}, /* 0x2465 */
            {8'h00}, /* 0x2464 */
            {8'h00}, /* 0x2463 */
            {8'h00}, /* 0x2462 */
            {8'h00}, /* 0x2461 */
            {8'h00}, /* 0x2460 */
            {8'h00}, /* 0x245f */
            {8'h00}, /* 0x245e */
            {8'h00}, /* 0x245d */
            {8'h00}, /* 0x245c */
            {8'h00}, /* 0x245b */
            {8'h00}, /* 0x245a */
            {8'h00}, /* 0x2459 */
            {8'h00}, /* 0x2458 */
            {8'h00}, /* 0x2457 */
            {8'h00}, /* 0x2456 */
            {8'h00}, /* 0x2455 */
            {8'h00}, /* 0x2454 */
            {8'h00}, /* 0x2453 */
            {8'h00}, /* 0x2452 */
            {8'h00}, /* 0x2451 */
            {8'h00}, /* 0x2450 */
            {8'h00}, /* 0x244f */
            {8'h00}, /* 0x244e */
            {8'h00}, /* 0x244d */
            {8'h00}, /* 0x244c */
            {8'h00}, /* 0x244b */
            {8'h00}, /* 0x244a */
            {8'h00}, /* 0x2449 */
            {8'h00}, /* 0x2448 */
            {8'h00}, /* 0x2447 */
            {8'h00}, /* 0x2446 */
            {8'h00}, /* 0x2445 */
            {8'h00}, /* 0x2444 */
            {8'h00}, /* 0x2443 */
            {8'h00}, /* 0x2442 */
            {8'h00}, /* 0x2441 */
            {8'h00}, /* 0x2440 */
            {8'h00}, /* 0x243f */
            {8'h00}, /* 0x243e */
            {8'h00}, /* 0x243d */
            {8'h00}, /* 0x243c */
            {8'h00}, /* 0x243b */
            {8'h00}, /* 0x243a */
            {8'h00}, /* 0x2439 */
            {8'h00}, /* 0x2438 */
            {8'h00}, /* 0x2437 */
            {8'h00}, /* 0x2436 */
            {8'h00}, /* 0x2435 */
            {8'h00}, /* 0x2434 */
            {8'h00}, /* 0x2433 */
            {8'h00}, /* 0x2432 */
            {8'h00}, /* 0x2431 */
            {8'h00}, /* 0x2430 */
            {8'h00}, /* 0x242f */
            {8'h00}, /* 0x242e */
            {8'h00}, /* 0x242d */
            {8'h00}, /* 0x242c */
            {8'h00}, /* 0x242b */
            {8'h00}, /* 0x242a */
            {8'h00}, /* 0x2429 */
            {8'h00}, /* 0x2428 */
            {8'h00}, /* 0x2427 */
            {8'h00}, /* 0x2426 */
            {8'h00}, /* 0x2425 */
            {8'h00}, /* 0x2424 */
            {8'h00}, /* 0x2423 */
            {8'h00}, /* 0x2422 */
            {8'h00}, /* 0x2421 */
            {8'h00}, /* 0x2420 */
            {8'h00}, /* 0x241f */
            {8'h00}, /* 0x241e */
            {8'h00}, /* 0x241d */
            {8'h00}, /* 0x241c */
            {8'h00}, /* 0x241b */
            {8'h00}, /* 0x241a */
            {8'h00}, /* 0x2419 */
            {8'h00}, /* 0x2418 */
            {8'h00}, /* 0x2417 */
            {8'h00}, /* 0x2416 */
            {8'h00}, /* 0x2415 */
            {8'h00}, /* 0x2414 */
            {8'h00}, /* 0x2413 */
            {8'h00}, /* 0x2412 */
            {8'h00}, /* 0x2411 */
            {8'h00}, /* 0x2410 */
            {8'h00}, /* 0x240f */
            {8'h00}, /* 0x240e */
            {8'h00}, /* 0x240d */
            {8'h00}, /* 0x240c */
            {8'h00}, /* 0x240b */
            {8'h00}, /* 0x240a */
            {8'h00}, /* 0x2409 */
            {8'h00}, /* 0x2408 */
            {8'h00}, /* 0x2407 */
            {8'h00}, /* 0x2406 */
            {8'h00}, /* 0x2405 */
            {8'h00}, /* 0x2404 */
            {8'h00}, /* 0x2403 */
            {8'h00}, /* 0x2402 */
            {8'h00}, /* 0x2401 */
            {8'h00}, /* 0x2400 */
            {8'h00}, /* 0x23ff */
            {8'h00}, /* 0x23fe */
            {8'h00}, /* 0x23fd */
            {8'h00}, /* 0x23fc */
            {8'h00}, /* 0x23fb */
            {8'h00}, /* 0x23fa */
            {8'h00}, /* 0x23f9 */
            {8'h00}, /* 0x23f8 */
            {8'h00}, /* 0x23f7 */
            {8'h00}, /* 0x23f6 */
            {8'h00}, /* 0x23f5 */
            {8'h00}, /* 0x23f4 */
            {8'h00}, /* 0x23f3 */
            {8'h00}, /* 0x23f2 */
            {8'h00}, /* 0x23f1 */
            {8'h00}, /* 0x23f0 */
            {8'h00}, /* 0x23ef */
            {8'h00}, /* 0x23ee */
            {8'h00}, /* 0x23ed */
            {8'h00}, /* 0x23ec */
            {8'h00}, /* 0x23eb */
            {8'h00}, /* 0x23ea */
            {8'h00}, /* 0x23e9 */
            {8'h00}, /* 0x23e8 */
            {8'h00}, /* 0x23e7 */
            {8'h00}, /* 0x23e6 */
            {8'h00}, /* 0x23e5 */
            {8'h00}, /* 0x23e4 */
            {8'h00}, /* 0x23e3 */
            {8'h00}, /* 0x23e2 */
            {8'h00}, /* 0x23e1 */
            {8'h00}, /* 0x23e0 */
            {8'h00}, /* 0x23df */
            {8'h00}, /* 0x23de */
            {8'h00}, /* 0x23dd */
            {8'h00}, /* 0x23dc */
            {8'h00}, /* 0x23db */
            {8'h00}, /* 0x23da */
            {8'h00}, /* 0x23d9 */
            {8'h00}, /* 0x23d8 */
            {8'h00}, /* 0x23d7 */
            {8'h00}, /* 0x23d6 */
            {8'h00}, /* 0x23d5 */
            {8'h00}, /* 0x23d4 */
            {8'h00}, /* 0x23d3 */
            {8'h00}, /* 0x23d2 */
            {8'h00}, /* 0x23d1 */
            {8'h00}, /* 0x23d0 */
            {8'h00}, /* 0x23cf */
            {8'h00}, /* 0x23ce */
            {8'h00}, /* 0x23cd */
            {8'h00}, /* 0x23cc */
            {8'h00}, /* 0x23cb */
            {8'h00}, /* 0x23ca */
            {8'h00}, /* 0x23c9 */
            {8'h00}, /* 0x23c8 */
            {8'h00}, /* 0x23c7 */
            {8'h00}, /* 0x23c6 */
            {8'h00}, /* 0x23c5 */
            {8'h00}, /* 0x23c4 */
            {8'h00}, /* 0x23c3 */
            {8'h00}, /* 0x23c2 */
            {8'h00}, /* 0x23c1 */
            {8'h00}, /* 0x23c0 */
            {8'h00}, /* 0x23bf */
            {8'h00}, /* 0x23be */
            {8'h00}, /* 0x23bd */
            {8'h00}, /* 0x23bc */
            {8'h00}, /* 0x23bb */
            {8'h00}, /* 0x23ba */
            {8'h00}, /* 0x23b9 */
            {8'h00}, /* 0x23b8 */
            {8'h00}, /* 0x23b7 */
            {8'h00}, /* 0x23b6 */
            {8'h00}, /* 0x23b5 */
            {8'h00}, /* 0x23b4 */
            {8'h00}, /* 0x23b3 */
            {8'h00}, /* 0x23b2 */
            {8'h00}, /* 0x23b1 */
            {8'h00}, /* 0x23b0 */
            {8'h00}, /* 0x23af */
            {8'h00}, /* 0x23ae */
            {8'h00}, /* 0x23ad */
            {8'h00}, /* 0x23ac */
            {8'h00}, /* 0x23ab */
            {8'h00}, /* 0x23aa */
            {8'h00}, /* 0x23a9 */
            {8'h00}, /* 0x23a8 */
            {8'h00}, /* 0x23a7 */
            {8'h00}, /* 0x23a6 */
            {8'h00}, /* 0x23a5 */
            {8'h00}, /* 0x23a4 */
            {8'h00}, /* 0x23a3 */
            {8'h00}, /* 0x23a2 */
            {8'h00}, /* 0x23a1 */
            {8'h00}, /* 0x23a0 */
            {8'h00}, /* 0x239f */
            {8'h00}, /* 0x239e */
            {8'h00}, /* 0x239d */
            {8'h00}, /* 0x239c */
            {8'h00}, /* 0x239b */
            {8'h00}, /* 0x239a */
            {8'h00}, /* 0x2399 */
            {8'h00}, /* 0x2398 */
            {8'h00}, /* 0x2397 */
            {8'h00}, /* 0x2396 */
            {8'h00}, /* 0x2395 */
            {8'h00}, /* 0x2394 */
            {8'h00}, /* 0x2393 */
            {8'h00}, /* 0x2392 */
            {8'h00}, /* 0x2391 */
            {8'h00}, /* 0x2390 */
            {8'h00}, /* 0x238f */
            {8'h00}, /* 0x238e */
            {8'h00}, /* 0x238d */
            {8'h00}, /* 0x238c */
            {8'h00}, /* 0x238b */
            {8'h00}, /* 0x238a */
            {8'h00}, /* 0x2389 */
            {8'h00}, /* 0x2388 */
            {8'h00}, /* 0x2387 */
            {8'h00}, /* 0x2386 */
            {8'h00}, /* 0x2385 */
            {8'h00}, /* 0x2384 */
            {8'h00}, /* 0x2383 */
            {8'h00}, /* 0x2382 */
            {8'h00}, /* 0x2381 */
            {8'h00}, /* 0x2380 */
            {8'h00}, /* 0x237f */
            {8'h00}, /* 0x237e */
            {8'h00}, /* 0x237d */
            {8'h00}, /* 0x237c */
            {8'h00}, /* 0x237b */
            {8'h00}, /* 0x237a */
            {8'h00}, /* 0x2379 */
            {8'h00}, /* 0x2378 */
            {8'h00}, /* 0x2377 */
            {8'h00}, /* 0x2376 */
            {8'h00}, /* 0x2375 */
            {8'h00}, /* 0x2374 */
            {8'h00}, /* 0x2373 */
            {8'h00}, /* 0x2372 */
            {8'h00}, /* 0x2371 */
            {8'h00}, /* 0x2370 */
            {8'h00}, /* 0x236f */
            {8'h00}, /* 0x236e */
            {8'h00}, /* 0x236d */
            {8'h00}, /* 0x236c */
            {8'h00}, /* 0x236b */
            {8'h00}, /* 0x236a */
            {8'h00}, /* 0x2369 */
            {8'h00}, /* 0x2368 */
            {8'h00}, /* 0x2367 */
            {8'h00}, /* 0x2366 */
            {8'h00}, /* 0x2365 */
            {8'h00}, /* 0x2364 */
            {8'h00}, /* 0x2363 */
            {8'h00}, /* 0x2362 */
            {8'h00}, /* 0x2361 */
            {8'h00}, /* 0x2360 */
            {8'h00}, /* 0x235f */
            {8'h00}, /* 0x235e */
            {8'h00}, /* 0x235d */
            {8'h00}, /* 0x235c */
            {8'h00}, /* 0x235b */
            {8'h00}, /* 0x235a */
            {8'h00}, /* 0x2359 */
            {8'h00}, /* 0x2358 */
            {8'h00}, /* 0x2357 */
            {8'h00}, /* 0x2356 */
            {8'h00}, /* 0x2355 */
            {8'h00}, /* 0x2354 */
            {8'h00}, /* 0x2353 */
            {8'h00}, /* 0x2352 */
            {8'h00}, /* 0x2351 */
            {8'h00}, /* 0x2350 */
            {8'h00}, /* 0x234f */
            {8'h00}, /* 0x234e */
            {8'h00}, /* 0x234d */
            {8'h00}, /* 0x234c */
            {8'h00}, /* 0x234b */
            {8'h00}, /* 0x234a */
            {8'h00}, /* 0x2349 */
            {8'h00}, /* 0x2348 */
            {8'h00}, /* 0x2347 */
            {8'h00}, /* 0x2346 */
            {8'h00}, /* 0x2345 */
            {8'h00}, /* 0x2344 */
            {8'h00}, /* 0x2343 */
            {8'h00}, /* 0x2342 */
            {8'h00}, /* 0x2341 */
            {8'h00}, /* 0x2340 */
            {8'h00}, /* 0x233f */
            {8'h00}, /* 0x233e */
            {8'h00}, /* 0x233d */
            {8'h00}, /* 0x233c */
            {8'h00}, /* 0x233b */
            {8'h00}, /* 0x233a */
            {8'h00}, /* 0x2339 */
            {8'h00}, /* 0x2338 */
            {8'h00}, /* 0x2337 */
            {8'h00}, /* 0x2336 */
            {8'h00}, /* 0x2335 */
            {8'h00}, /* 0x2334 */
            {8'h00}, /* 0x2333 */
            {8'h00}, /* 0x2332 */
            {8'h00}, /* 0x2331 */
            {8'h00}, /* 0x2330 */
            {8'h00}, /* 0x232f */
            {8'h00}, /* 0x232e */
            {8'h00}, /* 0x232d */
            {8'h00}, /* 0x232c */
            {8'h00}, /* 0x232b */
            {8'h00}, /* 0x232a */
            {8'h00}, /* 0x2329 */
            {8'h00}, /* 0x2328 */
            {8'h00}, /* 0x2327 */
            {8'h00}, /* 0x2326 */
            {8'h00}, /* 0x2325 */
            {8'h00}, /* 0x2324 */
            {8'h00}, /* 0x2323 */
            {8'h00}, /* 0x2322 */
            {8'h00}, /* 0x2321 */
            {8'h00}, /* 0x2320 */
            {8'h00}, /* 0x231f */
            {8'h00}, /* 0x231e */
            {8'h00}, /* 0x231d */
            {8'h00}, /* 0x231c */
            {8'h00}, /* 0x231b */
            {8'h00}, /* 0x231a */
            {8'h00}, /* 0x2319 */
            {8'h00}, /* 0x2318 */
            {8'h00}, /* 0x2317 */
            {8'h00}, /* 0x2316 */
            {8'h00}, /* 0x2315 */
            {8'h00}, /* 0x2314 */
            {8'h00}, /* 0x2313 */
            {8'h00}, /* 0x2312 */
            {8'h00}, /* 0x2311 */
            {8'h00}, /* 0x2310 */
            {8'h00}, /* 0x230f */
            {8'h00}, /* 0x230e */
            {8'h00}, /* 0x230d */
            {8'h00}, /* 0x230c */
            {8'h00}, /* 0x230b */
            {8'h00}, /* 0x230a */
            {8'h00}, /* 0x2309 */
            {8'h00}, /* 0x2308 */
            {8'h00}, /* 0x2307 */
            {8'h00}, /* 0x2306 */
            {8'h00}, /* 0x2305 */
            {8'h00}, /* 0x2304 */
            {8'h00}, /* 0x2303 */
            {8'h00}, /* 0x2302 */
            {8'h00}, /* 0x2301 */
            {8'h00}, /* 0x2300 */
            {8'h00}, /* 0x22ff */
            {8'h00}, /* 0x22fe */
            {8'h00}, /* 0x22fd */
            {8'h00}, /* 0x22fc */
            {8'h00}, /* 0x22fb */
            {8'h00}, /* 0x22fa */
            {8'h00}, /* 0x22f9 */
            {8'h00}, /* 0x22f8 */
            {8'h00}, /* 0x22f7 */
            {8'h00}, /* 0x22f6 */
            {8'h00}, /* 0x22f5 */
            {8'h00}, /* 0x22f4 */
            {8'h00}, /* 0x22f3 */
            {8'h00}, /* 0x22f2 */
            {8'h00}, /* 0x22f1 */
            {8'h00}, /* 0x22f0 */
            {8'h00}, /* 0x22ef */
            {8'h00}, /* 0x22ee */
            {8'h00}, /* 0x22ed */
            {8'h00}, /* 0x22ec */
            {8'h00}, /* 0x22eb */
            {8'h00}, /* 0x22ea */
            {8'h00}, /* 0x22e9 */
            {8'h00}, /* 0x22e8 */
            {8'h00}, /* 0x22e7 */
            {8'h00}, /* 0x22e6 */
            {8'h00}, /* 0x22e5 */
            {8'h00}, /* 0x22e4 */
            {8'h00}, /* 0x22e3 */
            {8'h00}, /* 0x22e2 */
            {8'h00}, /* 0x22e1 */
            {8'h00}, /* 0x22e0 */
            {8'h00}, /* 0x22df */
            {8'h00}, /* 0x22de */
            {8'h00}, /* 0x22dd */
            {8'h00}, /* 0x22dc */
            {8'h00}, /* 0x22db */
            {8'h00}, /* 0x22da */
            {8'h00}, /* 0x22d9 */
            {8'h00}, /* 0x22d8 */
            {8'h00}, /* 0x22d7 */
            {8'h00}, /* 0x22d6 */
            {8'h00}, /* 0x22d5 */
            {8'h00}, /* 0x22d4 */
            {8'h00}, /* 0x22d3 */
            {8'h00}, /* 0x22d2 */
            {8'h00}, /* 0x22d1 */
            {8'h00}, /* 0x22d0 */
            {8'h00}, /* 0x22cf */
            {8'h00}, /* 0x22ce */
            {8'h00}, /* 0x22cd */
            {8'h00}, /* 0x22cc */
            {8'h00}, /* 0x22cb */
            {8'h00}, /* 0x22ca */
            {8'h00}, /* 0x22c9 */
            {8'h00}, /* 0x22c8 */
            {8'h00}, /* 0x22c7 */
            {8'h00}, /* 0x22c6 */
            {8'h00}, /* 0x22c5 */
            {8'h00}, /* 0x22c4 */
            {8'h00}, /* 0x22c3 */
            {8'h00}, /* 0x22c2 */
            {8'h00}, /* 0x22c1 */
            {8'h00}, /* 0x22c0 */
            {8'h00}, /* 0x22bf */
            {8'h00}, /* 0x22be */
            {8'h00}, /* 0x22bd */
            {8'h00}, /* 0x22bc */
            {8'h00}, /* 0x22bb */
            {8'h00}, /* 0x22ba */
            {8'h00}, /* 0x22b9 */
            {8'h00}, /* 0x22b8 */
            {8'h00}, /* 0x22b7 */
            {8'h00}, /* 0x22b6 */
            {8'h00}, /* 0x22b5 */
            {8'h00}, /* 0x22b4 */
            {8'h00}, /* 0x22b3 */
            {8'h00}, /* 0x22b2 */
            {8'h00}, /* 0x22b1 */
            {8'h00}, /* 0x22b0 */
            {8'h00}, /* 0x22af */
            {8'h00}, /* 0x22ae */
            {8'h00}, /* 0x22ad */
            {8'h00}, /* 0x22ac */
            {8'h00}, /* 0x22ab */
            {8'h00}, /* 0x22aa */
            {8'h00}, /* 0x22a9 */
            {8'h00}, /* 0x22a8 */
            {8'h00}, /* 0x22a7 */
            {8'h00}, /* 0x22a6 */
            {8'h00}, /* 0x22a5 */
            {8'h00}, /* 0x22a4 */
            {8'h00}, /* 0x22a3 */
            {8'h00}, /* 0x22a2 */
            {8'h00}, /* 0x22a1 */
            {8'h00}, /* 0x22a0 */
            {8'h00}, /* 0x229f */
            {8'h00}, /* 0x229e */
            {8'h00}, /* 0x229d */
            {8'h00}, /* 0x229c */
            {8'h00}, /* 0x229b */
            {8'h00}, /* 0x229a */
            {8'h00}, /* 0x2299 */
            {8'h00}, /* 0x2298 */
            {8'h00}, /* 0x2297 */
            {8'h00}, /* 0x2296 */
            {8'h00}, /* 0x2295 */
            {8'h00}, /* 0x2294 */
            {8'h00}, /* 0x2293 */
            {8'h00}, /* 0x2292 */
            {8'h00}, /* 0x2291 */
            {8'h00}, /* 0x2290 */
            {8'h00}, /* 0x228f */
            {8'h00}, /* 0x228e */
            {8'h00}, /* 0x228d */
            {8'h00}, /* 0x228c */
            {8'h00}, /* 0x228b */
            {8'h00}, /* 0x228a */
            {8'h00}, /* 0x2289 */
            {8'h00}, /* 0x2288 */
            {8'h00}, /* 0x2287 */
            {8'h00}, /* 0x2286 */
            {8'h00}, /* 0x2285 */
            {8'h00}, /* 0x2284 */
            {8'h00}, /* 0x2283 */
            {8'h00}, /* 0x2282 */
            {8'h00}, /* 0x2281 */
            {8'h00}, /* 0x2280 */
            {8'h00}, /* 0x227f */
            {8'h00}, /* 0x227e */
            {8'h00}, /* 0x227d */
            {8'h00}, /* 0x227c */
            {8'h00}, /* 0x227b */
            {8'h00}, /* 0x227a */
            {8'h00}, /* 0x2279 */
            {8'h00}, /* 0x2278 */
            {8'h00}, /* 0x2277 */
            {8'h00}, /* 0x2276 */
            {8'h00}, /* 0x2275 */
            {8'h00}, /* 0x2274 */
            {8'h00}, /* 0x2273 */
            {8'h00}, /* 0x2272 */
            {8'h00}, /* 0x2271 */
            {8'h00}, /* 0x2270 */
            {8'h00}, /* 0x226f */
            {8'h00}, /* 0x226e */
            {8'h00}, /* 0x226d */
            {8'h00}, /* 0x226c */
            {8'h00}, /* 0x226b */
            {8'h00}, /* 0x226a */
            {8'h00}, /* 0x2269 */
            {8'h00}, /* 0x2268 */
            {8'h00}, /* 0x2267 */
            {8'h00}, /* 0x2266 */
            {8'h00}, /* 0x2265 */
            {8'h00}, /* 0x2264 */
            {8'h00}, /* 0x2263 */
            {8'h00}, /* 0x2262 */
            {8'h00}, /* 0x2261 */
            {8'h00}, /* 0x2260 */
            {8'h00}, /* 0x225f */
            {8'h00}, /* 0x225e */
            {8'h00}, /* 0x225d */
            {8'h00}, /* 0x225c */
            {8'h00}, /* 0x225b */
            {8'h00}, /* 0x225a */
            {8'h00}, /* 0x2259 */
            {8'h00}, /* 0x2258 */
            {8'h00}, /* 0x2257 */
            {8'h00}, /* 0x2256 */
            {8'h00}, /* 0x2255 */
            {8'h00}, /* 0x2254 */
            {8'h00}, /* 0x2253 */
            {8'h00}, /* 0x2252 */
            {8'h00}, /* 0x2251 */
            {8'h00}, /* 0x2250 */
            {8'h00}, /* 0x224f */
            {8'h00}, /* 0x224e */
            {8'h00}, /* 0x224d */
            {8'h00}, /* 0x224c */
            {8'h00}, /* 0x224b */
            {8'h00}, /* 0x224a */
            {8'h00}, /* 0x2249 */
            {8'h00}, /* 0x2248 */
            {8'h00}, /* 0x2247 */
            {8'h00}, /* 0x2246 */
            {8'h00}, /* 0x2245 */
            {8'h00}, /* 0x2244 */
            {8'h00}, /* 0x2243 */
            {8'h00}, /* 0x2242 */
            {8'h00}, /* 0x2241 */
            {8'h00}, /* 0x2240 */
            {8'h00}, /* 0x223f */
            {8'h00}, /* 0x223e */
            {8'h00}, /* 0x223d */
            {8'h00}, /* 0x223c */
            {8'h00}, /* 0x223b */
            {8'h00}, /* 0x223a */
            {8'h00}, /* 0x2239 */
            {8'h00}, /* 0x2238 */
            {8'h00}, /* 0x2237 */
            {8'h00}, /* 0x2236 */
            {8'h00}, /* 0x2235 */
            {8'h00}, /* 0x2234 */
            {8'h00}, /* 0x2233 */
            {8'h00}, /* 0x2232 */
            {8'h00}, /* 0x2231 */
            {8'h00}, /* 0x2230 */
            {8'h00}, /* 0x222f */
            {8'h00}, /* 0x222e */
            {8'h00}, /* 0x222d */
            {8'h00}, /* 0x222c */
            {8'h00}, /* 0x222b */
            {8'h00}, /* 0x222a */
            {8'h00}, /* 0x2229 */
            {8'h00}, /* 0x2228 */
            {8'h00}, /* 0x2227 */
            {8'h00}, /* 0x2226 */
            {8'h00}, /* 0x2225 */
            {8'h00}, /* 0x2224 */
            {8'h00}, /* 0x2223 */
            {8'h00}, /* 0x2222 */
            {8'h00}, /* 0x2221 */
            {8'h00}, /* 0x2220 */
            {8'h00}, /* 0x221f */
            {8'h00}, /* 0x221e */
            {8'h00}, /* 0x221d */
            {8'h00}, /* 0x221c */
            {8'h00}, /* 0x221b */
            {8'h00}, /* 0x221a */
            {8'h00}, /* 0x2219 */
            {8'h00}, /* 0x2218 */
            {8'h00}, /* 0x2217 */
            {8'h00}, /* 0x2216 */
            {8'h00}, /* 0x2215 */
            {8'h00}, /* 0x2214 */
            {8'h00}, /* 0x2213 */
            {8'h00}, /* 0x2212 */
            {8'h00}, /* 0x2211 */
            {8'h00}, /* 0x2210 */
            {8'h00}, /* 0x220f */
            {8'h00}, /* 0x220e */
            {8'h00}, /* 0x220d */
            {8'h00}, /* 0x220c */
            {8'h00}, /* 0x220b */
            {8'h00}, /* 0x220a */
            {8'h00}, /* 0x2209 */
            {8'h00}, /* 0x2208 */
            {8'h00}, /* 0x2207 */
            {8'h00}, /* 0x2206 */
            {8'h00}, /* 0x2205 */
            {8'h00}, /* 0x2204 */
            {8'h00}, /* 0x2203 */
            {8'h00}, /* 0x2202 */
            {8'h00}, /* 0x2201 */
            {8'h00}, /* 0x2200 */
            {8'h00}, /* 0x21ff */
            {8'h00}, /* 0x21fe */
            {8'h00}, /* 0x21fd */
            {8'h00}, /* 0x21fc */
            {8'h00}, /* 0x21fb */
            {8'h00}, /* 0x21fa */
            {8'h00}, /* 0x21f9 */
            {8'h00}, /* 0x21f8 */
            {8'h00}, /* 0x21f7 */
            {8'h00}, /* 0x21f6 */
            {8'h00}, /* 0x21f5 */
            {8'h00}, /* 0x21f4 */
            {8'h00}, /* 0x21f3 */
            {8'h00}, /* 0x21f2 */
            {8'h00}, /* 0x21f1 */
            {8'h00}, /* 0x21f0 */
            {8'h00}, /* 0x21ef */
            {8'h00}, /* 0x21ee */
            {8'h00}, /* 0x21ed */
            {8'h00}, /* 0x21ec */
            {8'h00}, /* 0x21eb */
            {8'h00}, /* 0x21ea */
            {8'h00}, /* 0x21e9 */
            {8'h00}, /* 0x21e8 */
            {8'h00}, /* 0x21e7 */
            {8'h00}, /* 0x21e6 */
            {8'h00}, /* 0x21e5 */
            {8'h00}, /* 0x21e4 */
            {8'h00}, /* 0x21e3 */
            {8'h00}, /* 0x21e2 */
            {8'h00}, /* 0x21e1 */
            {8'h00}, /* 0x21e0 */
            {8'h00}, /* 0x21df */
            {8'h00}, /* 0x21de */
            {8'h00}, /* 0x21dd */
            {8'h00}, /* 0x21dc */
            {8'h00}, /* 0x21db */
            {8'h00}, /* 0x21da */
            {8'h00}, /* 0x21d9 */
            {8'h00}, /* 0x21d8 */
            {8'h00}, /* 0x21d7 */
            {8'h00}, /* 0x21d6 */
            {8'h00}, /* 0x21d5 */
            {8'h00}, /* 0x21d4 */
            {8'h00}, /* 0x21d3 */
            {8'h00}, /* 0x21d2 */
            {8'h00}, /* 0x21d1 */
            {8'h00}, /* 0x21d0 */
            {8'h00}, /* 0x21cf */
            {8'h00}, /* 0x21ce */
            {8'h00}, /* 0x21cd */
            {8'h00}, /* 0x21cc */
            {8'h00}, /* 0x21cb */
            {8'h00}, /* 0x21ca */
            {8'h00}, /* 0x21c9 */
            {8'h00}, /* 0x21c8 */
            {8'h00}, /* 0x21c7 */
            {8'h00}, /* 0x21c6 */
            {8'h00}, /* 0x21c5 */
            {8'h00}, /* 0x21c4 */
            {8'h00}, /* 0x21c3 */
            {8'h00}, /* 0x21c2 */
            {8'h00}, /* 0x21c1 */
            {8'h00}, /* 0x21c0 */
            {8'h00}, /* 0x21bf */
            {8'h00}, /* 0x21be */
            {8'h00}, /* 0x21bd */
            {8'h00}, /* 0x21bc */
            {8'h00}, /* 0x21bb */
            {8'h00}, /* 0x21ba */
            {8'h00}, /* 0x21b9 */
            {8'h00}, /* 0x21b8 */
            {8'h00}, /* 0x21b7 */
            {8'h00}, /* 0x21b6 */
            {8'h00}, /* 0x21b5 */
            {8'h00}, /* 0x21b4 */
            {8'h00}, /* 0x21b3 */
            {8'h00}, /* 0x21b2 */
            {8'h00}, /* 0x21b1 */
            {8'h00}, /* 0x21b0 */
            {8'h00}, /* 0x21af */
            {8'h00}, /* 0x21ae */
            {8'h00}, /* 0x21ad */
            {8'h00}, /* 0x21ac */
            {8'h00}, /* 0x21ab */
            {8'h00}, /* 0x21aa */
            {8'h00}, /* 0x21a9 */
            {8'h00}, /* 0x21a8 */
            {8'h00}, /* 0x21a7 */
            {8'h00}, /* 0x21a6 */
            {8'h00}, /* 0x21a5 */
            {8'h00}, /* 0x21a4 */
            {8'h00}, /* 0x21a3 */
            {8'h00}, /* 0x21a2 */
            {8'h00}, /* 0x21a1 */
            {8'h00}, /* 0x21a0 */
            {8'h00}, /* 0x219f */
            {8'h00}, /* 0x219e */
            {8'h00}, /* 0x219d */
            {8'h00}, /* 0x219c */
            {8'h00}, /* 0x219b */
            {8'h00}, /* 0x219a */
            {8'h00}, /* 0x2199 */
            {8'h00}, /* 0x2198 */
            {8'h00}, /* 0x2197 */
            {8'h00}, /* 0x2196 */
            {8'h00}, /* 0x2195 */
            {8'h00}, /* 0x2194 */
            {8'h00}, /* 0x2193 */
            {8'h00}, /* 0x2192 */
            {8'h00}, /* 0x2191 */
            {8'h00}, /* 0x2190 */
            {8'h00}, /* 0x218f */
            {8'h00}, /* 0x218e */
            {8'h00}, /* 0x218d */
            {8'h00}, /* 0x218c */
            {8'h00}, /* 0x218b */
            {8'h00}, /* 0x218a */
            {8'h00}, /* 0x2189 */
            {8'h00}, /* 0x2188 */
            {8'h00}, /* 0x2187 */
            {8'h00}, /* 0x2186 */
            {8'h00}, /* 0x2185 */
            {8'h00}, /* 0x2184 */
            {8'h00}, /* 0x2183 */
            {8'h00}, /* 0x2182 */
            {8'h00}, /* 0x2181 */
            {8'h00}, /* 0x2180 */
            {8'h00}, /* 0x217f */
            {8'h00}, /* 0x217e */
            {8'h00}, /* 0x217d */
            {8'h00}, /* 0x217c */
            {8'h00}, /* 0x217b */
            {8'h00}, /* 0x217a */
            {8'h00}, /* 0x2179 */
            {8'h00}, /* 0x2178 */
            {8'h00}, /* 0x2177 */
            {8'h00}, /* 0x2176 */
            {8'h00}, /* 0x2175 */
            {8'h00}, /* 0x2174 */
            {8'h00}, /* 0x2173 */
            {8'h00}, /* 0x2172 */
            {8'h00}, /* 0x2171 */
            {8'h00}, /* 0x2170 */
            {8'h00}, /* 0x216f */
            {8'h00}, /* 0x216e */
            {8'h00}, /* 0x216d */
            {8'h00}, /* 0x216c */
            {8'h00}, /* 0x216b */
            {8'h00}, /* 0x216a */
            {8'h00}, /* 0x2169 */
            {8'h00}, /* 0x2168 */
            {8'h00}, /* 0x2167 */
            {8'h00}, /* 0x2166 */
            {8'h00}, /* 0x2165 */
            {8'h00}, /* 0x2164 */
            {8'h00}, /* 0x2163 */
            {8'h00}, /* 0x2162 */
            {8'h00}, /* 0x2161 */
            {8'h00}, /* 0x2160 */
            {8'h00}, /* 0x215f */
            {8'h00}, /* 0x215e */
            {8'h00}, /* 0x215d */
            {8'h00}, /* 0x215c */
            {8'h00}, /* 0x215b */
            {8'h00}, /* 0x215a */
            {8'h00}, /* 0x2159 */
            {8'h00}, /* 0x2158 */
            {8'h00}, /* 0x2157 */
            {8'h00}, /* 0x2156 */
            {8'h00}, /* 0x2155 */
            {8'h00}, /* 0x2154 */
            {8'h00}, /* 0x2153 */
            {8'h00}, /* 0x2152 */
            {8'h00}, /* 0x2151 */
            {8'h00}, /* 0x2150 */
            {8'h00}, /* 0x214f */
            {8'h00}, /* 0x214e */
            {8'h00}, /* 0x214d */
            {8'h00}, /* 0x214c */
            {8'h00}, /* 0x214b */
            {8'h00}, /* 0x214a */
            {8'h00}, /* 0x2149 */
            {8'h00}, /* 0x2148 */
            {8'h00}, /* 0x2147 */
            {8'h00}, /* 0x2146 */
            {8'h00}, /* 0x2145 */
            {8'h00}, /* 0x2144 */
            {8'h00}, /* 0x2143 */
            {8'h00}, /* 0x2142 */
            {8'h00}, /* 0x2141 */
            {8'h00}, /* 0x2140 */
            {8'h00}, /* 0x213f */
            {8'h00}, /* 0x213e */
            {8'h00}, /* 0x213d */
            {8'h00}, /* 0x213c */
            {8'h00}, /* 0x213b */
            {8'h00}, /* 0x213a */
            {8'h00}, /* 0x2139 */
            {8'h00}, /* 0x2138 */
            {8'h00}, /* 0x2137 */
            {8'h00}, /* 0x2136 */
            {8'h00}, /* 0x2135 */
            {8'h00}, /* 0x2134 */
            {8'h00}, /* 0x2133 */
            {8'h00}, /* 0x2132 */
            {8'h00}, /* 0x2131 */
            {8'h00}, /* 0x2130 */
            {8'h00}, /* 0x212f */
            {8'h00}, /* 0x212e */
            {8'h00}, /* 0x212d */
            {8'h00}, /* 0x212c */
            {8'h00}, /* 0x212b */
            {8'h00}, /* 0x212a */
            {8'h00}, /* 0x2129 */
            {8'h00}, /* 0x2128 */
            {8'h00}, /* 0x2127 */
            {8'h00}, /* 0x2126 */
            {8'h00}, /* 0x2125 */
            {8'h00}, /* 0x2124 */
            {8'h00}, /* 0x2123 */
            {8'h00}, /* 0x2122 */
            {8'h00}, /* 0x2121 */
            {8'h00}, /* 0x2120 */
            {8'h00}, /* 0x211f */
            {8'h00}, /* 0x211e */
            {8'h00}, /* 0x211d */
            {8'h00}, /* 0x211c */
            {8'h00}, /* 0x211b */
            {8'h00}, /* 0x211a */
            {8'h00}, /* 0x2119 */
            {8'h00}, /* 0x2118 */
            {8'h00}, /* 0x2117 */
            {8'h00}, /* 0x2116 */
            {8'h00}, /* 0x2115 */
            {8'h00}, /* 0x2114 */
            {8'h00}, /* 0x2113 */
            {8'h00}, /* 0x2112 */
            {8'h00}, /* 0x2111 */
            {8'h00}, /* 0x2110 */
            {8'h00}, /* 0x210f */
            {8'h00}, /* 0x210e */
            {8'h00}, /* 0x210d */
            {8'h00}, /* 0x210c */
            {8'h00}, /* 0x210b */
            {8'h00}, /* 0x210a */
            {8'h00}, /* 0x2109 */
            {8'h00}, /* 0x2108 */
            {8'h00}, /* 0x2107 */
            {8'h00}, /* 0x2106 */
            {8'h00}, /* 0x2105 */
            {8'h00}, /* 0x2104 */
            {8'h00}, /* 0x2103 */
            {8'h00}, /* 0x2102 */
            {8'h00}, /* 0x2101 */
            {8'h00}, /* 0x2100 */
            {8'h00}, /* 0x20ff */
            {8'h00}, /* 0x20fe */
            {8'h00}, /* 0x20fd */
            {8'h00}, /* 0x20fc */
            {8'h00}, /* 0x20fb */
            {8'h00}, /* 0x20fa */
            {8'h00}, /* 0x20f9 */
            {8'h00}, /* 0x20f8 */
            {8'h00}, /* 0x20f7 */
            {8'h00}, /* 0x20f6 */
            {8'h00}, /* 0x20f5 */
            {8'h00}, /* 0x20f4 */
            {8'h00}, /* 0x20f3 */
            {8'h00}, /* 0x20f2 */
            {8'h00}, /* 0x20f1 */
            {8'h00}, /* 0x20f0 */
            {8'h00}, /* 0x20ef */
            {8'h00}, /* 0x20ee */
            {8'h00}, /* 0x20ed */
            {8'h00}, /* 0x20ec */
            {8'h00}, /* 0x20eb */
            {8'h00}, /* 0x20ea */
            {8'h00}, /* 0x20e9 */
            {8'h00}, /* 0x20e8 */
            {8'h00}, /* 0x20e7 */
            {8'h00}, /* 0x20e6 */
            {8'h00}, /* 0x20e5 */
            {8'h00}, /* 0x20e4 */
            {8'h00}, /* 0x20e3 */
            {8'h00}, /* 0x20e2 */
            {8'h00}, /* 0x20e1 */
            {8'h00}, /* 0x20e0 */
            {8'h00}, /* 0x20df */
            {8'h00}, /* 0x20de */
            {8'h00}, /* 0x20dd */
            {8'h00}, /* 0x20dc */
            {8'h00}, /* 0x20db */
            {8'h00}, /* 0x20da */
            {8'h00}, /* 0x20d9 */
            {8'h00}, /* 0x20d8 */
            {8'h00}, /* 0x20d7 */
            {8'h00}, /* 0x20d6 */
            {8'h00}, /* 0x20d5 */
            {8'h00}, /* 0x20d4 */
            {8'h00}, /* 0x20d3 */
            {8'h00}, /* 0x20d2 */
            {8'h00}, /* 0x20d1 */
            {8'h00}, /* 0x20d0 */
            {8'h00}, /* 0x20cf */
            {8'h00}, /* 0x20ce */
            {8'h00}, /* 0x20cd */
            {8'h00}, /* 0x20cc */
            {8'h00}, /* 0x20cb */
            {8'h00}, /* 0x20ca */
            {8'h00}, /* 0x20c9 */
            {8'h00}, /* 0x20c8 */
            {8'h00}, /* 0x20c7 */
            {8'h00}, /* 0x20c6 */
            {8'h00}, /* 0x20c5 */
            {8'h00}, /* 0x20c4 */
            {8'h00}, /* 0x20c3 */
            {8'h00}, /* 0x20c2 */
            {8'h00}, /* 0x20c1 */
            {8'h00}, /* 0x20c0 */
            {8'h00}, /* 0x20bf */
            {8'h00}, /* 0x20be */
            {8'h00}, /* 0x20bd */
            {8'h00}, /* 0x20bc */
            {8'h00}, /* 0x20bb */
            {8'h00}, /* 0x20ba */
            {8'h00}, /* 0x20b9 */
            {8'h00}, /* 0x20b8 */
            {8'h00}, /* 0x20b7 */
            {8'h00}, /* 0x20b6 */
            {8'h00}, /* 0x20b5 */
            {8'h00}, /* 0x20b4 */
            {8'h00}, /* 0x20b3 */
            {8'h00}, /* 0x20b2 */
            {8'h00}, /* 0x20b1 */
            {8'h00}, /* 0x20b0 */
            {8'h00}, /* 0x20af */
            {8'h00}, /* 0x20ae */
            {8'h00}, /* 0x20ad */
            {8'h00}, /* 0x20ac */
            {8'h00}, /* 0x20ab */
            {8'h00}, /* 0x20aa */
            {8'h00}, /* 0x20a9 */
            {8'h00}, /* 0x20a8 */
            {8'h00}, /* 0x20a7 */
            {8'h00}, /* 0x20a6 */
            {8'h00}, /* 0x20a5 */
            {8'h00}, /* 0x20a4 */
            {8'h00}, /* 0x20a3 */
            {8'h00}, /* 0x20a2 */
            {8'h00}, /* 0x20a1 */
            {8'h00}, /* 0x20a0 */
            {8'h00}, /* 0x209f */
            {8'h00}, /* 0x209e */
            {8'h00}, /* 0x209d */
            {8'h00}, /* 0x209c */
            {8'h00}, /* 0x209b */
            {8'h00}, /* 0x209a */
            {8'h00}, /* 0x2099 */
            {8'h00}, /* 0x2098 */
            {8'h00}, /* 0x2097 */
            {8'h00}, /* 0x2096 */
            {8'h00}, /* 0x2095 */
            {8'h00}, /* 0x2094 */
            {8'h00}, /* 0x2093 */
            {8'h00}, /* 0x2092 */
            {8'h00}, /* 0x2091 */
            {8'h00}, /* 0x2090 */
            {8'h00}, /* 0x208f */
            {8'h00}, /* 0x208e */
            {8'h00}, /* 0x208d */
            {8'h00}, /* 0x208c */
            {8'h00}, /* 0x208b */
            {8'h00}, /* 0x208a */
            {8'h00}, /* 0x2089 */
            {8'h00}, /* 0x2088 */
            {8'h00}, /* 0x2087 */
            {8'h00}, /* 0x2086 */
            {8'h00}, /* 0x2085 */
            {8'h00}, /* 0x2084 */
            {8'h00}, /* 0x2083 */
            {8'h00}, /* 0x2082 */
            {8'h00}, /* 0x2081 */
            {8'h00}, /* 0x2080 */
            {8'h00}, /* 0x207f */
            {8'h00}, /* 0x207e */
            {8'h00}, /* 0x207d */
            {8'h00}, /* 0x207c */
            {8'h00}, /* 0x207b */
            {8'h00}, /* 0x207a */
            {8'h00}, /* 0x2079 */
            {8'h00}, /* 0x2078 */
            {8'h00}, /* 0x2077 */
            {8'h00}, /* 0x2076 */
            {8'h00}, /* 0x2075 */
            {8'h00}, /* 0x2074 */
            {8'h00}, /* 0x2073 */
            {8'h00}, /* 0x2072 */
            {8'h00}, /* 0x2071 */
            {8'h00}, /* 0x2070 */
            {8'h00}, /* 0x206f */
            {8'h00}, /* 0x206e */
            {8'h00}, /* 0x206d */
            {8'h00}, /* 0x206c */
            {8'h00}, /* 0x206b */
            {8'h00}, /* 0x206a */
            {8'h00}, /* 0x2069 */
            {8'h00}, /* 0x2068 */
            {8'h00}, /* 0x2067 */
            {8'h00}, /* 0x2066 */
            {8'h00}, /* 0x2065 */
            {8'h00}, /* 0x2064 */
            {8'h00}, /* 0x2063 */
            {8'h00}, /* 0x2062 */
            {8'h00}, /* 0x2061 */
            {8'h00}, /* 0x2060 */
            {8'h00}, /* 0x205f */
            {8'h00}, /* 0x205e */
            {8'h00}, /* 0x205d */
            {8'h00}, /* 0x205c */
            {8'h00}, /* 0x205b */
            {8'h00}, /* 0x205a */
            {8'h00}, /* 0x2059 */
            {8'h00}, /* 0x2058 */
            {8'h00}, /* 0x2057 */
            {8'h00}, /* 0x2056 */
            {8'h00}, /* 0x2055 */
            {8'h00}, /* 0x2054 */
            {8'h00}, /* 0x2053 */
            {8'h00}, /* 0x2052 */
            {8'h00}, /* 0x2051 */
            {8'h00}, /* 0x2050 */
            {8'h00}, /* 0x204f */
            {8'h00}, /* 0x204e */
            {8'h00}, /* 0x204d */
            {8'h00}, /* 0x204c */
            {8'h00}, /* 0x204b */
            {8'h00}, /* 0x204a */
            {8'h00}, /* 0x2049 */
            {8'h00}, /* 0x2048 */
            {8'h00}, /* 0x2047 */
            {8'h00}, /* 0x2046 */
            {8'h00}, /* 0x2045 */
            {8'h00}, /* 0x2044 */
            {8'h00}, /* 0x2043 */
            {8'h00}, /* 0x2042 */
            {8'h00}, /* 0x2041 */
            {8'h00}, /* 0x2040 */
            {8'h00}, /* 0x203f */
            {8'h00}, /* 0x203e */
            {8'h00}, /* 0x203d */
            {8'h00}, /* 0x203c */
            {8'h00}, /* 0x203b */
            {8'h00}, /* 0x203a */
            {8'h00}, /* 0x2039 */
            {8'h00}, /* 0x2038 */
            {8'h00}, /* 0x2037 */
            {8'h00}, /* 0x2036 */
            {8'h00}, /* 0x2035 */
            {8'h00}, /* 0x2034 */
            {8'h00}, /* 0x2033 */
            {8'h00}, /* 0x2032 */
            {8'h00}, /* 0x2031 */
            {8'h00}, /* 0x2030 */
            {8'h00}, /* 0x202f */
            {8'h00}, /* 0x202e */
            {8'h00}, /* 0x202d */
            {8'h00}, /* 0x202c */
            {8'h00}, /* 0x202b */
            {8'h00}, /* 0x202a */
            {8'h00}, /* 0x2029 */
            {8'h00}, /* 0x2028 */
            {8'h00}, /* 0x2027 */
            {8'h00}, /* 0x2026 */
            {8'h00}, /* 0x2025 */
            {8'h00}, /* 0x2024 */
            {8'h00}, /* 0x2023 */
            {8'h00}, /* 0x2022 */
            {8'h00}, /* 0x2021 */
            {8'h00}, /* 0x2020 */
            {8'h00}, /* 0x201f */
            {8'h00}, /* 0x201e */
            {8'h00}, /* 0x201d */
            {8'h00}, /* 0x201c */
            {8'h00}, /* 0x201b */
            {8'h00}, /* 0x201a */
            {8'h00}, /* 0x2019 */
            {8'h00}, /* 0x2018 */
            {8'h00}, /* 0x2017 */
            {8'h00}, /* 0x2016 */
            {8'h00}, /* 0x2015 */
            {8'h00}, /* 0x2014 */
            {8'h00}, /* 0x2013 */
            {8'h00}, /* 0x2012 */
            {8'h00}, /* 0x2011 */
            {8'h00}, /* 0x2010 */
            {8'h00}, /* 0x200f */
            {8'h00}, /* 0x200e */
            {8'h00}, /* 0x200d */
            {8'h00}, /* 0x200c */
            {8'h00}, /* 0x200b */
            {8'h00}, /* 0x200a */
            {8'h00}, /* 0x2009 */
            {8'h00}, /* 0x2008 */
            {8'h00}, /* 0x2007 */
            {8'h00}, /* 0x2006 */
            {8'h00}, /* 0x2005 */
            {8'h00}, /* 0x2004 */
            {8'h00}, /* 0x2003 */
            {8'h00}, /* 0x2002 */
            {8'h00}, /* 0x2001 */
            {8'h00}, /* 0x2000 */
            {8'h00}, /* 0x1fff */
            {8'h00}, /* 0x1ffe */
            {8'h00}, /* 0x1ffd */
            {8'h00}, /* 0x1ffc */
            {8'h00}, /* 0x1ffb */
            {8'h00}, /* 0x1ffa */
            {8'h00}, /* 0x1ff9 */
            {8'h00}, /* 0x1ff8 */
            {8'h00}, /* 0x1ff7 */
            {8'h00}, /* 0x1ff6 */
            {8'h00}, /* 0x1ff5 */
            {8'h00}, /* 0x1ff4 */
            {8'h00}, /* 0x1ff3 */
            {8'h00}, /* 0x1ff2 */
            {8'h00}, /* 0x1ff1 */
            {8'h00}, /* 0x1ff0 */
            {8'h00}, /* 0x1fef */
            {8'h00}, /* 0x1fee */
            {8'h00}, /* 0x1fed */
            {8'h00}, /* 0x1fec */
            {8'h00}, /* 0x1feb */
            {8'h00}, /* 0x1fea */
            {8'h00}, /* 0x1fe9 */
            {8'h00}, /* 0x1fe8 */
            {8'h00}, /* 0x1fe7 */
            {8'h00}, /* 0x1fe6 */
            {8'h00}, /* 0x1fe5 */
            {8'h00}, /* 0x1fe4 */
            {8'h00}, /* 0x1fe3 */
            {8'h00}, /* 0x1fe2 */
            {8'h00}, /* 0x1fe1 */
            {8'h00}, /* 0x1fe0 */
            {8'h00}, /* 0x1fdf */
            {8'h00}, /* 0x1fde */
            {8'h00}, /* 0x1fdd */
            {8'h00}, /* 0x1fdc */
            {8'h00}, /* 0x1fdb */
            {8'h00}, /* 0x1fda */
            {8'h00}, /* 0x1fd9 */
            {8'h00}, /* 0x1fd8 */
            {8'h00}, /* 0x1fd7 */
            {8'h00}, /* 0x1fd6 */
            {8'h00}, /* 0x1fd5 */
            {8'h00}, /* 0x1fd4 */
            {8'h00}, /* 0x1fd3 */
            {8'h00}, /* 0x1fd2 */
            {8'h00}, /* 0x1fd1 */
            {8'h00}, /* 0x1fd0 */
            {8'h00}, /* 0x1fcf */
            {8'h00}, /* 0x1fce */
            {8'h00}, /* 0x1fcd */
            {8'h00}, /* 0x1fcc */
            {8'h00}, /* 0x1fcb */
            {8'h00}, /* 0x1fca */
            {8'h00}, /* 0x1fc9 */
            {8'h00}, /* 0x1fc8 */
            {8'h00}, /* 0x1fc7 */
            {8'h00}, /* 0x1fc6 */
            {8'h00}, /* 0x1fc5 */
            {8'h00}, /* 0x1fc4 */
            {8'h00}, /* 0x1fc3 */
            {8'h00}, /* 0x1fc2 */
            {8'h00}, /* 0x1fc1 */
            {8'h00}, /* 0x1fc0 */
            {8'h00}, /* 0x1fbf */
            {8'h00}, /* 0x1fbe */
            {8'h00}, /* 0x1fbd */
            {8'h00}, /* 0x1fbc */
            {8'h00}, /* 0x1fbb */
            {8'h00}, /* 0x1fba */
            {8'h00}, /* 0x1fb9 */
            {8'h00}, /* 0x1fb8 */
            {8'h00}, /* 0x1fb7 */
            {8'h00}, /* 0x1fb6 */
            {8'h00}, /* 0x1fb5 */
            {8'h00}, /* 0x1fb4 */
            {8'h00}, /* 0x1fb3 */
            {8'h00}, /* 0x1fb2 */
            {8'h00}, /* 0x1fb1 */
            {8'h00}, /* 0x1fb0 */
            {8'h00}, /* 0x1faf */
            {8'h00}, /* 0x1fae */
            {8'h00}, /* 0x1fad */
            {8'h00}, /* 0x1fac */
            {8'h00}, /* 0x1fab */
            {8'h00}, /* 0x1faa */
            {8'h00}, /* 0x1fa9 */
            {8'h00}, /* 0x1fa8 */
            {8'h00}, /* 0x1fa7 */
            {8'h00}, /* 0x1fa6 */
            {8'h00}, /* 0x1fa5 */
            {8'h00}, /* 0x1fa4 */
            {8'h00}, /* 0x1fa3 */
            {8'h00}, /* 0x1fa2 */
            {8'h00}, /* 0x1fa1 */
            {8'h00}, /* 0x1fa0 */
            {8'h00}, /* 0x1f9f */
            {8'h00}, /* 0x1f9e */
            {8'h00}, /* 0x1f9d */
            {8'h00}, /* 0x1f9c */
            {8'h00}, /* 0x1f9b */
            {8'h00}, /* 0x1f9a */
            {8'h00}, /* 0x1f99 */
            {8'h00}, /* 0x1f98 */
            {8'h00}, /* 0x1f97 */
            {8'h00}, /* 0x1f96 */
            {8'h00}, /* 0x1f95 */
            {8'h00}, /* 0x1f94 */
            {8'h00}, /* 0x1f93 */
            {8'h00}, /* 0x1f92 */
            {8'h00}, /* 0x1f91 */
            {8'h00}, /* 0x1f90 */
            {8'h00}, /* 0x1f8f */
            {8'h00}, /* 0x1f8e */
            {8'h00}, /* 0x1f8d */
            {8'h00}, /* 0x1f8c */
            {8'h00}, /* 0x1f8b */
            {8'h00}, /* 0x1f8a */
            {8'h00}, /* 0x1f89 */
            {8'h00}, /* 0x1f88 */
            {8'h00}, /* 0x1f87 */
            {8'h00}, /* 0x1f86 */
            {8'h00}, /* 0x1f85 */
            {8'h00}, /* 0x1f84 */
            {8'h00}, /* 0x1f83 */
            {8'h00}, /* 0x1f82 */
            {8'h00}, /* 0x1f81 */
            {8'h00}, /* 0x1f80 */
            {8'h00}, /* 0x1f7f */
            {8'h00}, /* 0x1f7e */
            {8'h00}, /* 0x1f7d */
            {8'h00}, /* 0x1f7c */
            {8'h00}, /* 0x1f7b */
            {8'h00}, /* 0x1f7a */
            {8'h00}, /* 0x1f79 */
            {8'h00}, /* 0x1f78 */
            {8'h00}, /* 0x1f77 */
            {8'h00}, /* 0x1f76 */
            {8'h00}, /* 0x1f75 */
            {8'h00}, /* 0x1f74 */
            {8'h00}, /* 0x1f73 */
            {8'h00}, /* 0x1f72 */
            {8'h00}, /* 0x1f71 */
            {8'h00}, /* 0x1f70 */
            {8'h00}, /* 0x1f6f */
            {8'h00}, /* 0x1f6e */
            {8'h00}, /* 0x1f6d */
            {8'h00}, /* 0x1f6c */
            {8'h00}, /* 0x1f6b */
            {8'h00}, /* 0x1f6a */
            {8'h00}, /* 0x1f69 */
            {8'h00}, /* 0x1f68 */
            {8'h00}, /* 0x1f67 */
            {8'h00}, /* 0x1f66 */
            {8'h00}, /* 0x1f65 */
            {8'h00}, /* 0x1f64 */
            {8'h00}, /* 0x1f63 */
            {8'h00}, /* 0x1f62 */
            {8'h00}, /* 0x1f61 */
            {8'h00}, /* 0x1f60 */
            {8'h00}, /* 0x1f5f */
            {8'h00}, /* 0x1f5e */
            {8'h00}, /* 0x1f5d */
            {8'h00}, /* 0x1f5c */
            {8'h00}, /* 0x1f5b */
            {8'h00}, /* 0x1f5a */
            {8'h00}, /* 0x1f59 */
            {8'h00}, /* 0x1f58 */
            {8'h00}, /* 0x1f57 */
            {8'h00}, /* 0x1f56 */
            {8'h00}, /* 0x1f55 */
            {8'h00}, /* 0x1f54 */
            {8'h00}, /* 0x1f53 */
            {8'h00}, /* 0x1f52 */
            {8'h00}, /* 0x1f51 */
            {8'h00}, /* 0x1f50 */
            {8'h00}, /* 0x1f4f */
            {8'h00}, /* 0x1f4e */
            {8'h00}, /* 0x1f4d */
            {8'h00}, /* 0x1f4c */
            {8'h00}, /* 0x1f4b */
            {8'h00}, /* 0x1f4a */
            {8'h00}, /* 0x1f49 */
            {8'h00}, /* 0x1f48 */
            {8'h00}, /* 0x1f47 */
            {8'h00}, /* 0x1f46 */
            {8'h00}, /* 0x1f45 */
            {8'h00}, /* 0x1f44 */
            {8'h00}, /* 0x1f43 */
            {8'h00}, /* 0x1f42 */
            {8'h00}, /* 0x1f41 */
            {8'h00}, /* 0x1f40 */
            {8'h00}, /* 0x1f3f */
            {8'h00}, /* 0x1f3e */
            {8'h00}, /* 0x1f3d */
            {8'h00}, /* 0x1f3c */
            {8'h00}, /* 0x1f3b */
            {8'h00}, /* 0x1f3a */
            {8'h00}, /* 0x1f39 */
            {8'h00}, /* 0x1f38 */
            {8'h00}, /* 0x1f37 */
            {8'h00}, /* 0x1f36 */
            {8'h00}, /* 0x1f35 */
            {8'h00}, /* 0x1f34 */
            {8'h00}, /* 0x1f33 */
            {8'h00}, /* 0x1f32 */
            {8'h00}, /* 0x1f31 */
            {8'h00}, /* 0x1f30 */
            {8'h00}, /* 0x1f2f */
            {8'h00}, /* 0x1f2e */
            {8'h00}, /* 0x1f2d */
            {8'h00}, /* 0x1f2c */
            {8'h00}, /* 0x1f2b */
            {8'h00}, /* 0x1f2a */
            {8'h00}, /* 0x1f29 */
            {8'h00}, /* 0x1f28 */
            {8'h00}, /* 0x1f27 */
            {8'h00}, /* 0x1f26 */
            {8'h00}, /* 0x1f25 */
            {8'h00}, /* 0x1f24 */
            {8'h00}, /* 0x1f23 */
            {8'h00}, /* 0x1f22 */
            {8'h00}, /* 0x1f21 */
            {8'h00}, /* 0x1f20 */
            {8'h00}, /* 0x1f1f */
            {8'h00}, /* 0x1f1e */
            {8'h00}, /* 0x1f1d */
            {8'h00}, /* 0x1f1c */
            {8'h00}, /* 0x1f1b */
            {8'h00}, /* 0x1f1a */
            {8'h00}, /* 0x1f19 */
            {8'h00}, /* 0x1f18 */
            {8'h00}, /* 0x1f17 */
            {8'h00}, /* 0x1f16 */
            {8'h00}, /* 0x1f15 */
            {8'h00}, /* 0x1f14 */
            {8'h00}, /* 0x1f13 */
            {8'h00}, /* 0x1f12 */
            {8'h00}, /* 0x1f11 */
            {8'h00}, /* 0x1f10 */
            {8'h00}, /* 0x1f0f */
            {8'h00}, /* 0x1f0e */
            {8'h00}, /* 0x1f0d */
            {8'h00}, /* 0x1f0c */
            {8'h00}, /* 0x1f0b */
            {8'h00}, /* 0x1f0a */
            {8'h00}, /* 0x1f09 */
            {8'h00}, /* 0x1f08 */
            {8'h00}, /* 0x1f07 */
            {8'h00}, /* 0x1f06 */
            {8'h00}, /* 0x1f05 */
            {8'h00}, /* 0x1f04 */
            {8'h00}, /* 0x1f03 */
            {8'h00}, /* 0x1f02 */
            {8'h00}, /* 0x1f01 */
            {8'h00}, /* 0x1f00 */
            {8'h00}, /* 0x1eff */
            {8'h00}, /* 0x1efe */
            {8'h00}, /* 0x1efd */
            {8'h00}, /* 0x1efc */
            {8'h00}, /* 0x1efb */
            {8'h00}, /* 0x1efa */
            {8'h00}, /* 0x1ef9 */
            {8'h00}, /* 0x1ef8 */
            {8'h00}, /* 0x1ef7 */
            {8'h00}, /* 0x1ef6 */
            {8'h00}, /* 0x1ef5 */
            {8'h00}, /* 0x1ef4 */
            {8'h00}, /* 0x1ef3 */
            {8'h00}, /* 0x1ef2 */
            {8'h00}, /* 0x1ef1 */
            {8'h00}, /* 0x1ef0 */
            {8'h00}, /* 0x1eef */
            {8'h00}, /* 0x1eee */
            {8'h00}, /* 0x1eed */
            {8'h00}, /* 0x1eec */
            {8'h00}, /* 0x1eeb */
            {8'h00}, /* 0x1eea */
            {8'h00}, /* 0x1ee9 */
            {8'h00}, /* 0x1ee8 */
            {8'h00}, /* 0x1ee7 */
            {8'h00}, /* 0x1ee6 */
            {8'h00}, /* 0x1ee5 */
            {8'h00}, /* 0x1ee4 */
            {8'h00}, /* 0x1ee3 */
            {8'h00}, /* 0x1ee2 */
            {8'h00}, /* 0x1ee1 */
            {8'h00}, /* 0x1ee0 */
            {8'h00}, /* 0x1edf */
            {8'h00}, /* 0x1ede */
            {8'h00}, /* 0x1edd */
            {8'h00}, /* 0x1edc */
            {8'h00}, /* 0x1edb */
            {8'h00}, /* 0x1eda */
            {8'h00}, /* 0x1ed9 */
            {8'h00}, /* 0x1ed8 */
            {8'h00}, /* 0x1ed7 */
            {8'h00}, /* 0x1ed6 */
            {8'h00}, /* 0x1ed5 */
            {8'h00}, /* 0x1ed4 */
            {8'h00}, /* 0x1ed3 */
            {8'h00}, /* 0x1ed2 */
            {8'h00}, /* 0x1ed1 */
            {8'h00}, /* 0x1ed0 */
            {8'h00}, /* 0x1ecf */
            {8'h00}, /* 0x1ece */
            {8'h00}, /* 0x1ecd */
            {8'h00}, /* 0x1ecc */
            {8'h00}, /* 0x1ecb */
            {8'h00}, /* 0x1eca */
            {8'h00}, /* 0x1ec9 */
            {8'h00}, /* 0x1ec8 */
            {8'h00}, /* 0x1ec7 */
            {8'h00}, /* 0x1ec6 */
            {8'h00}, /* 0x1ec5 */
            {8'h00}, /* 0x1ec4 */
            {8'h00}, /* 0x1ec3 */
            {8'h00}, /* 0x1ec2 */
            {8'h00}, /* 0x1ec1 */
            {8'h00}, /* 0x1ec0 */
            {8'h00}, /* 0x1ebf */
            {8'h00}, /* 0x1ebe */
            {8'h00}, /* 0x1ebd */
            {8'h00}, /* 0x1ebc */
            {8'h00}, /* 0x1ebb */
            {8'h00}, /* 0x1eba */
            {8'h00}, /* 0x1eb9 */
            {8'h00}, /* 0x1eb8 */
            {8'h00}, /* 0x1eb7 */
            {8'h00}, /* 0x1eb6 */
            {8'h00}, /* 0x1eb5 */
            {8'h00}, /* 0x1eb4 */
            {8'h00}, /* 0x1eb3 */
            {8'h00}, /* 0x1eb2 */
            {8'h00}, /* 0x1eb1 */
            {8'h00}, /* 0x1eb0 */
            {8'h00}, /* 0x1eaf */
            {8'h00}, /* 0x1eae */
            {8'h00}, /* 0x1ead */
            {8'h00}, /* 0x1eac */
            {8'h00}, /* 0x1eab */
            {8'h00}, /* 0x1eaa */
            {8'h00}, /* 0x1ea9 */
            {8'h00}, /* 0x1ea8 */
            {8'h00}, /* 0x1ea7 */
            {8'h00}, /* 0x1ea6 */
            {8'h00}, /* 0x1ea5 */
            {8'h00}, /* 0x1ea4 */
            {8'h00}, /* 0x1ea3 */
            {8'h00}, /* 0x1ea2 */
            {8'h00}, /* 0x1ea1 */
            {8'h00}, /* 0x1ea0 */
            {8'h00}, /* 0x1e9f */
            {8'h00}, /* 0x1e9e */
            {8'h00}, /* 0x1e9d */
            {8'h00}, /* 0x1e9c */
            {8'h00}, /* 0x1e9b */
            {8'h00}, /* 0x1e9a */
            {8'h00}, /* 0x1e99 */
            {8'h00}, /* 0x1e98 */
            {8'h00}, /* 0x1e97 */
            {8'h00}, /* 0x1e96 */
            {8'h00}, /* 0x1e95 */
            {8'h00}, /* 0x1e94 */
            {8'h00}, /* 0x1e93 */
            {8'h00}, /* 0x1e92 */
            {8'h00}, /* 0x1e91 */
            {8'h00}, /* 0x1e90 */
            {8'h00}, /* 0x1e8f */
            {8'h00}, /* 0x1e8e */
            {8'h00}, /* 0x1e8d */
            {8'h00}, /* 0x1e8c */
            {8'h00}, /* 0x1e8b */
            {8'h00}, /* 0x1e8a */
            {8'h00}, /* 0x1e89 */
            {8'h00}, /* 0x1e88 */
            {8'h00}, /* 0x1e87 */
            {8'h00}, /* 0x1e86 */
            {8'h00}, /* 0x1e85 */
            {8'h00}, /* 0x1e84 */
            {8'h00}, /* 0x1e83 */
            {8'h00}, /* 0x1e82 */
            {8'h00}, /* 0x1e81 */
            {8'h00}, /* 0x1e80 */
            {8'h00}, /* 0x1e7f */
            {8'h00}, /* 0x1e7e */
            {8'h00}, /* 0x1e7d */
            {8'h00}, /* 0x1e7c */
            {8'h00}, /* 0x1e7b */
            {8'h00}, /* 0x1e7a */
            {8'h00}, /* 0x1e79 */
            {8'h00}, /* 0x1e78 */
            {8'h00}, /* 0x1e77 */
            {8'h00}, /* 0x1e76 */
            {8'h00}, /* 0x1e75 */
            {8'h00}, /* 0x1e74 */
            {8'h00}, /* 0x1e73 */
            {8'h00}, /* 0x1e72 */
            {8'h00}, /* 0x1e71 */
            {8'h00}, /* 0x1e70 */
            {8'h00}, /* 0x1e6f */
            {8'h00}, /* 0x1e6e */
            {8'h00}, /* 0x1e6d */
            {8'h00}, /* 0x1e6c */
            {8'h00}, /* 0x1e6b */
            {8'h00}, /* 0x1e6a */
            {8'h00}, /* 0x1e69 */
            {8'h00}, /* 0x1e68 */
            {8'h00}, /* 0x1e67 */
            {8'h00}, /* 0x1e66 */
            {8'h00}, /* 0x1e65 */
            {8'h00}, /* 0x1e64 */
            {8'h00}, /* 0x1e63 */
            {8'h00}, /* 0x1e62 */
            {8'h00}, /* 0x1e61 */
            {8'h00}, /* 0x1e60 */
            {8'h00}, /* 0x1e5f */
            {8'h00}, /* 0x1e5e */
            {8'h00}, /* 0x1e5d */
            {8'h00}, /* 0x1e5c */
            {8'h00}, /* 0x1e5b */
            {8'h00}, /* 0x1e5a */
            {8'h00}, /* 0x1e59 */
            {8'h00}, /* 0x1e58 */
            {8'h00}, /* 0x1e57 */
            {8'h00}, /* 0x1e56 */
            {8'h00}, /* 0x1e55 */
            {8'h00}, /* 0x1e54 */
            {8'h00}, /* 0x1e53 */
            {8'h00}, /* 0x1e52 */
            {8'h00}, /* 0x1e51 */
            {8'h00}, /* 0x1e50 */
            {8'h00}, /* 0x1e4f */
            {8'h00}, /* 0x1e4e */
            {8'h00}, /* 0x1e4d */
            {8'h00}, /* 0x1e4c */
            {8'h00}, /* 0x1e4b */
            {8'h00}, /* 0x1e4a */
            {8'h00}, /* 0x1e49 */
            {8'h00}, /* 0x1e48 */
            {8'h00}, /* 0x1e47 */
            {8'h00}, /* 0x1e46 */
            {8'h00}, /* 0x1e45 */
            {8'h00}, /* 0x1e44 */
            {8'h00}, /* 0x1e43 */
            {8'h00}, /* 0x1e42 */
            {8'h00}, /* 0x1e41 */
            {8'h00}, /* 0x1e40 */
            {8'h00}, /* 0x1e3f */
            {8'h00}, /* 0x1e3e */
            {8'h00}, /* 0x1e3d */
            {8'h00}, /* 0x1e3c */
            {8'h00}, /* 0x1e3b */
            {8'h00}, /* 0x1e3a */
            {8'h00}, /* 0x1e39 */
            {8'h00}, /* 0x1e38 */
            {8'h00}, /* 0x1e37 */
            {8'h00}, /* 0x1e36 */
            {8'h00}, /* 0x1e35 */
            {8'h00}, /* 0x1e34 */
            {8'h00}, /* 0x1e33 */
            {8'h00}, /* 0x1e32 */
            {8'h00}, /* 0x1e31 */
            {8'h00}, /* 0x1e30 */
            {8'h00}, /* 0x1e2f */
            {8'h00}, /* 0x1e2e */
            {8'h00}, /* 0x1e2d */
            {8'h00}, /* 0x1e2c */
            {8'h00}, /* 0x1e2b */
            {8'h00}, /* 0x1e2a */
            {8'h00}, /* 0x1e29 */
            {8'h00}, /* 0x1e28 */
            {8'h00}, /* 0x1e27 */
            {8'h00}, /* 0x1e26 */
            {8'h00}, /* 0x1e25 */
            {8'h00}, /* 0x1e24 */
            {8'h00}, /* 0x1e23 */
            {8'h00}, /* 0x1e22 */
            {8'h00}, /* 0x1e21 */
            {8'h00}, /* 0x1e20 */
            {8'h00}, /* 0x1e1f */
            {8'h00}, /* 0x1e1e */
            {8'h00}, /* 0x1e1d */
            {8'h00}, /* 0x1e1c */
            {8'h00}, /* 0x1e1b */
            {8'h00}, /* 0x1e1a */
            {8'h00}, /* 0x1e19 */
            {8'h00}, /* 0x1e18 */
            {8'h00}, /* 0x1e17 */
            {8'h00}, /* 0x1e16 */
            {8'h00}, /* 0x1e15 */
            {8'h00}, /* 0x1e14 */
            {8'h00}, /* 0x1e13 */
            {8'h00}, /* 0x1e12 */
            {8'h00}, /* 0x1e11 */
            {8'h00}, /* 0x1e10 */
            {8'h00}, /* 0x1e0f */
            {8'h00}, /* 0x1e0e */
            {8'h00}, /* 0x1e0d */
            {8'h00}, /* 0x1e0c */
            {8'h00}, /* 0x1e0b */
            {8'h00}, /* 0x1e0a */
            {8'h00}, /* 0x1e09 */
            {8'h00}, /* 0x1e08 */
            {8'h00}, /* 0x1e07 */
            {8'h00}, /* 0x1e06 */
            {8'h00}, /* 0x1e05 */
            {8'h00}, /* 0x1e04 */
            {8'h00}, /* 0x1e03 */
            {8'h00}, /* 0x1e02 */
            {8'h00}, /* 0x1e01 */
            {8'h00}, /* 0x1e00 */
            {8'h00}, /* 0x1dff */
            {8'h00}, /* 0x1dfe */
            {8'h00}, /* 0x1dfd */
            {8'h00}, /* 0x1dfc */
            {8'h00}, /* 0x1dfb */
            {8'h00}, /* 0x1dfa */
            {8'h00}, /* 0x1df9 */
            {8'h00}, /* 0x1df8 */
            {8'h00}, /* 0x1df7 */
            {8'h00}, /* 0x1df6 */
            {8'h00}, /* 0x1df5 */
            {8'h00}, /* 0x1df4 */
            {8'h00}, /* 0x1df3 */
            {8'h00}, /* 0x1df2 */
            {8'h00}, /* 0x1df1 */
            {8'h00}, /* 0x1df0 */
            {8'h00}, /* 0x1def */
            {8'h00}, /* 0x1dee */
            {8'h00}, /* 0x1ded */
            {8'h00}, /* 0x1dec */
            {8'h00}, /* 0x1deb */
            {8'h00}, /* 0x1dea */
            {8'h00}, /* 0x1de9 */
            {8'h00}, /* 0x1de8 */
            {8'h00}, /* 0x1de7 */
            {8'h00}, /* 0x1de6 */
            {8'h00}, /* 0x1de5 */
            {8'h00}, /* 0x1de4 */
            {8'h00}, /* 0x1de3 */
            {8'h00}, /* 0x1de2 */
            {8'h00}, /* 0x1de1 */
            {8'h00}, /* 0x1de0 */
            {8'h00}, /* 0x1ddf */
            {8'h00}, /* 0x1dde */
            {8'h00}, /* 0x1ddd */
            {8'h00}, /* 0x1ddc */
            {8'h00}, /* 0x1ddb */
            {8'h00}, /* 0x1dda */
            {8'h00}, /* 0x1dd9 */
            {8'h00}, /* 0x1dd8 */
            {8'h00}, /* 0x1dd7 */
            {8'h00}, /* 0x1dd6 */
            {8'h00}, /* 0x1dd5 */
            {8'h00}, /* 0x1dd4 */
            {8'h00}, /* 0x1dd3 */
            {8'h00}, /* 0x1dd2 */
            {8'h00}, /* 0x1dd1 */
            {8'h00}, /* 0x1dd0 */
            {8'h00}, /* 0x1dcf */
            {8'h00}, /* 0x1dce */
            {8'h00}, /* 0x1dcd */
            {8'h00}, /* 0x1dcc */
            {8'h00}, /* 0x1dcb */
            {8'h00}, /* 0x1dca */
            {8'h00}, /* 0x1dc9 */
            {8'h00}, /* 0x1dc8 */
            {8'h00}, /* 0x1dc7 */
            {8'h00}, /* 0x1dc6 */
            {8'h00}, /* 0x1dc5 */
            {8'h00}, /* 0x1dc4 */
            {8'h00}, /* 0x1dc3 */
            {8'h00}, /* 0x1dc2 */
            {8'h00}, /* 0x1dc1 */
            {8'h00}, /* 0x1dc0 */
            {8'h00}, /* 0x1dbf */
            {8'h00}, /* 0x1dbe */
            {8'h00}, /* 0x1dbd */
            {8'h00}, /* 0x1dbc */
            {8'h00}, /* 0x1dbb */
            {8'h00}, /* 0x1dba */
            {8'h00}, /* 0x1db9 */
            {8'h00}, /* 0x1db8 */
            {8'h00}, /* 0x1db7 */
            {8'h00}, /* 0x1db6 */
            {8'h00}, /* 0x1db5 */
            {8'h00}, /* 0x1db4 */
            {8'h00}, /* 0x1db3 */
            {8'h00}, /* 0x1db2 */
            {8'h00}, /* 0x1db1 */
            {8'h00}, /* 0x1db0 */
            {8'h00}, /* 0x1daf */
            {8'h00}, /* 0x1dae */
            {8'h00}, /* 0x1dad */
            {8'h00}, /* 0x1dac */
            {8'h00}, /* 0x1dab */
            {8'h00}, /* 0x1daa */
            {8'h00}, /* 0x1da9 */
            {8'h00}, /* 0x1da8 */
            {8'h00}, /* 0x1da7 */
            {8'h00}, /* 0x1da6 */
            {8'h00}, /* 0x1da5 */
            {8'h00}, /* 0x1da4 */
            {8'h00}, /* 0x1da3 */
            {8'h00}, /* 0x1da2 */
            {8'h00}, /* 0x1da1 */
            {8'h00}, /* 0x1da0 */
            {8'h00}, /* 0x1d9f */
            {8'h00}, /* 0x1d9e */
            {8'h00}, /* 0x1d9d */
            {8'h00}, /* 0x1d9c */
            {8'h00}, /* 0x1d9b */
            {8'h00}, /* 0x1d9a */
            {8'h00}, /* 0x1d99 */
            {8'h00}, /* 0x1d98 */
            {8'h00}, /* 0x1d97 */
            {8'h00}, /* 0x1d96 */
            {8'h00}, /* 0x1d95 */
            {8'h00}, /* 0x1d94 */
            {8'h00}, /* 0x1d93 */
            {8'h00}, /* 0x1d92 */
            {8'h00}, /* 0x1d91 */
            {8'h00}, /* 0x1d90 */
            {8'h00}, /* 0x1d8f */
            {8'h00}, /* 0x1d8e */
            {8'h00}, /* 0x1d8d */
            {8'h00}, /* 0x1d8c */
            {8'h00}, /* 0x1d8b */
            {8'h00}, /* 0x1d8a */
            {8'h00}, /* 0x1d89 */
            {8'h00}, /* 0x1d88 */
            {8'h00}, /* 0x1d87 */
            {8'h00}, /* 0x1d86 */
            {8'h00}, /* 0x1d85 */
            {8'h00}, /* 0x1d84 */
            {8'h00}, /* 0x1d83 */
            {8'h00}, /* 0x1d82 */
            {8'h00}, /* 0x1d81 */
            {8'h00}, /* 0x1d80 */
            {8'h00}, /* 0x1d7f */
            {8'h00}, /* 0x1d7e */
            {8'h00}, /* 0x1d7d */
            {8'h00}, /* 0x1d7c */
            {8'h00}, /* 0x1d7b */
            {8'h00}, /* 0x1d7a */
            {8'h00}, /* 0x1d79 */
            {8'h00}, /* 0x1d78 */
            {8'h00}, /* 0x1d77 */
            {8'h00}, /* 0x1d76 */
            {8'h00}, /* 0x1d75 */
            {8'h00}, /* 0x1d74 */
            {8'h00}, /* 0x1d73 */
            {8'h00}, /* 0x1d72 */
            {8'h00}, /* 0x1d71 */
            {8'h00}, /* 0x1d70 */
            {8'h00}, /* 0x1d6f */
            {8'h00}, /* 0x1d6e */
            {8'h00}, /* 0x1d6d */
            {8'h00}, /* 0x1d6c */
            {8'h00}, /* 0x1d6b */
            {8'h00}, /* 0x1d6a */
            {8'h00}, /* 0x1d69 */
            {8'h00}, /* 0x1d68 */
            {8'h00}, /* 0x1d67 */
            {8'h00}, /* 0x1d66 */
            {8'h00}, /* 0x1d65 */
            {8'h00}, /* 0x1d64 */
            {8'h00}, /* 0x1d63 */
            {8'h00}, /* 0x1d62 */
            {8'h00}, /* 0x1d61 */
            {8'h00}, /* 0x1d60 */
            {8'h00}, /* 0x1d5f */
            {8'h00}, /* 0x1d5e */
            {8'h00}, /* 0x1d5d */
            {8'h00}, /* 0x1d5c */
            {8'h00}, /* 0x1d5b */
            {8'h00}, /* 0x1d5a */
            {8'h00}, /* 0x1d59 */
            {8'h00}, /* 0x1d58 */
            {8'h00}, /* 0x1d57 */
            {8'h00}, /* 0x1d56 */
            {8'h00}, /* 0x1d55 */
            {8'h00}, /* 0x1d54 */
            {8'h00}, /* 0x1d53 */
            {8'h00}, /* 0x1d52 */
            {8'h00}, /* 0x1d51 */
            {8'h00}, /* 0x1d50 */
            {8'h00}, /* 0x1d4f */
            {8'h00}, /* 0x1d4e */
            {8'h00}, /* 0x1d4d */
            {8'h00}, /* 0x1d4c */
            {8'h00}, /* 0x1d4b */
            {8'h00}, /* 0x1d4a */
            {8'h00}, /* 0x1d49 */
            {8'h00}, /* 0x1d48 */
            {8'h00}, /* 0x1d47 */
            {8'h00}, /* 0x1d46 */
            {8'h00}, /* 0x1d45 */
            {8'h00}, /* 0x1d44 */
            {8'h00}, /* 0x1d43 */
            {8'h00}, /* 0x1d42 */
            {8'h00}, /* 0x1d41 */
            {8'h00}, /* 0x1d40 */
            {8'h00}, /* 0x1d3f */
            {8'h00}, /* 0x1d3e */
            {8'h00}, /* 0x1d3d */
            {8'h00}, /* 0x1d3c */
            {8'h00}, /* 0x1d3b */
            {8'h00}, /* 0x1d3a */
            {8'h00}, /* 0x1d39 */
            {8'h00}, /* 0x1d38 */
            {8'h00}, /* 0x1d37 */
            {8'h00}, /* 0x1d36 */
            {8'h00}, /* 0x1d35 */
            {8'h00}, /* 0x1d34 */
            {8'h00}, /* 0x1d33 */
            {8'h00}, /* 0x1d32 */
            {8'h00}, /* 0x1d31 */
            {8'h00}, /* 0x1d30 */
            {8'h00}, /* 0x1d2f */
            {8'h00}, /* 0x1d2e */
            {8'h00}, /* 0x1d2d */
            {8'h00}, /* 0x1d2c */
            {8'h00}, /* 0x1d2b */
            {8'h00}, /* 0x1d2a */
            {8'h00}, /* 0x1d29 */
            {8'h00}, /* 0x1d28 */
            {8'h00}, /* 0x1d27 */
            {8'h00}, /* 0x1d26 */
            {8'h00}, /* 0x1d25 */
            {8'h00}, /* 0x1d24 */
            {8'h00}, /* 0x1d23 */
            {8'h00}, /* 0x1d22 */
            {8'h00}, /* 0x1d21 */
            {8'h00}, /* 0x1d20 */
            {8'h00}, /* 0x1d1f */
            {8'h00}, /* 0x1d1e */
            {8'h00}, /* 0x1d1d */
            {8'h00}, /* 0x1d1c */
            {8'h00}, /* 0x1d1b */
            {8'h00}, /* 0x1d1a */
            {8'h00}, /* 0x1d19 */
            {8'h00}, /* 0x1d18 */
            {8'h00}, /* 0x1d17 */
            {8'h00}, /* 0x1d16 */
            {8'h00}, /* 0x1d15 */
            {8'h00}, /* 0x1d14 */
            {8'h00}, /* 0x1d13 */
            {8'h00}, /* 0x1d12 */
            {8'h00}, /* 0x1d11 */
            {8'h00}, /* 0x1d10 */
            {8'h00}, /* 0x1d0f */
            {8'h00}, /* 0x1d0e */
            {8'h00}, /* 0x1d0d */
            {8'h00}, /* 0x1d0c */
            {8'h00}, /* 0x1d0b */
            {8'h00}, /* 0x1d0a */
            {8'h00}, /* 0x1d09 */
            {8'h00}, /* 0x1d08 */
            {8'h00}, /* 0x1d07 */
            {8'h00}, /* 0x1d06 */
            {8'h00}, /* 0x1d05 */
            {8'h00}, /* 0x1d04 */
            {8'h00}, /* 0x1d03 */
            {8'h00}, /* 0x1d02 */
            {8'h00}, /* 0x1d01 */
            {8'h00}, /* 0x1d00 */
            {8'h00}, /* 0x1cff */
            {8'h00}, /* 0x1cfe */
            {8'h00}, /* 0x1cfd */
            {8'h00}, /* 0x1cfc */
            {8'h00}, /* 0x1cfb */
            {8'h00}, /* 0x1cfa */
            {8'h00}, /* 0x1cf9 */
            {8'h00}, /* 0x1cf8 */
            {8'h00}, /* 0x1cf7 */
            {8'h00}, /* 0x1cf6 */
            {8'h00}, /* 0x1cf5 */
            {8'h00}, /* 0x1cf4 */
            {8'h00}, /* 0x1cf3 */
            {8'h00}, /* 0x1cf2 */
            {8'h00}, /* 0x1cf1 */
            {8'h00}, /* 0x1cf0 */
            {8'h00}, /* 0x1cef */
            {8'h00}, /* 0x1cee */
            {8'h00}, /* 0x1ced */
            {8'h00}, /* 0x1cec */
            {8'h00}, /* 0x1ceb */
            {8'h00}, /* 0x1cea */
            {8'h00}, /* 0x1ce9 */
            {8'h00}, /* 0x1ce8 */
            {8'h00}, /* 0x1ce7 */
            {8'h00}, /* 0x1ce6 */
            {8'h00}, /* 0x1ce5 */
            {8'h00}, /* 0x1ce4 */
            {8'h00}, /* 0x1ce3 */
            {8'h00}, /* 0x1ce2 */
            {8'h00}, /* 0x1ce1 */
            {8'h00}, /* 0x1ce0 */
            {8'h00}, /* 0x1cdf */
            {8'h00}, /* 0x1cde */
            {8'h00}, /* 0x1cdd */
            {8'h00}, /* 0x1cdc */
            {8'h00}, /* 0x1cdb */
            {8'h00}, /* 0x1cda */
            {8'h00}, /* 0x1cd9 */
            {8'h00}, /* 0x1cd8 */
            {8'h00}, /* 0x1cd7 */
            {8'h00}, /* 0x1cd6 */
            {8'h00}, /* 0x1cd5 */
            {8'h00}, /* 0x1cd4 */
            {8'h00}, /* 0x1cd3 */
            {8'h00}, /* 0x1cd2 */
            {8'h00}, /* 0x1cd1 */
            {8'h00}, /* 0x1cd0 */
            {8'h00}, /* 0x1ccf */
            {8'h00}, /* 0x1cce */
            {8'h00}, /* 0x1ccd */
            {8'h00}, /* 0x1ccc */
            {8'h00}, /* 0x1ccb */
            {8'h00}, /* 0x1cca */
            {8'h00}, /* 0x1cc9 */
            {8'h00}, /* 0x1cc8 */
            {8'h00}, /* 0x1cc7 */
            {8'h00}, /* 0x1cc6 */
            {8'h00}, /* 0x1cc5 */
            {8'h00}, /* 0x1cc4 */
            {8'h00}, /* 0x1cc3 */
            {8'h00}, /* 0x1cc2 */
            {8'h00}, /* 0x1cc1 */
            {8'h00}, /* 0x1cc0 */
            {8'h00}, /* 0x1cbf */
            {8'h00}, /* 0x1cbe */
            {8'h00}, /* 0x1cbd */
            {8'h00}, /* 0x1cbc */
            {8'h00}, /* 0x1cbb */
            {8'h00}, /* 0x1cba */
            {8'h00}, /* 0x1cb9 */
            {8'h00}, /* 0x1cb8 */
            {8'h00}, /* 0x1cb7 */
            {8'h00}, /* 0x1cb6 */
            {8'h00}, /* 0x1cb5 */
            {8'h00}, /* 0x1cb4 */
            {8'h00}, /* 0x1cb3 */
            {8'h00}, /* 0x1cb2 */
            {8'h00}, /* 0x1cb1 */
            {8'h00}, /* 0x1cb0 */
            {8'h00}, /* 0x1caf */
            {8'h00}, /* 0x1cae */
            {8'h00}, /* 0x1cad */
            {8'h00}, /* 0x1cac */
            {8'h00}, /* 0x1cab */
            {8'h00}, /* 0x1caa */
            {8'h00}, /* 0x1ca9 */
            {8'h00}, /* 0x1ca8 */
            {8'h00}, /* 0x1ca7 */
            {8'h00}, /* 0x1ca6 */
            {8'h00}, /* 0x1ca5 */
            {8'h00}, /* 0x1ca4 */
            {8'h00}, /* 0x1ca3 */
            {8'h00}, /* 0x1ca2 */
            {8'h00}, /* 0x1ca1 */
            {8'h00}, /* 0x1ca0 */
            {8'h00}, /* 0x1c9f */
            {8'h00}, /* 0x1c9e */
            {8'h00}, /* 0x1c9d */
            {8'h00}, /* 0x1c9c */
            {8'h00}, /* 0x1c9b */
            {8'h00}, /* 0x1c9a */
            {8'h00}, /* 0x1c99 */
            {8'h00}, /* 0x1c98 */
            {8'h00}, /* 0x1c97 */
            {8'h00}, /* 0x1c96 */
            {8'h00}, /* 0x1c95 */
            {8'h00}, /* 0x1c94 */
            {8'h00}, /* 0x1c93 */
            {8'h00}, /* 0x1c92 */
            {8'h00}, /* 0x1c91 */
            {8'h00}, /* 0x1c90 */
            {8'h00}, /* 0x1c8f */
            {8'h00}, /* 0x1c8e */
            {8'h00}, /* 0x1c8d */
            {8'h00}, /* 0x1c8c */
            {8'h00}, /* 0x1c8b */
            {8'h00}, /* 0x1c8a */
            {8'h00}, /* 0x1c89 */
            {8'h00}, /* 0x1c88 */
            {8'h00}, /* 0x1c87 */
            {8'h00}, /* 0x1c86 */
            {8'h00}, /* 0x1c85 */
            {8'h00}, /* 0x1c84 */
            {8'h00}, /* 0x1c83 */
            {8'h00}, /* 0x1c82 */
            {8'h00}, /* 0x1c81 */
            {8'h00}, /* 0x1c80 */
            {8'h00}, /* 0x1c7f */
            {8'h00}, /* 0x1c7e */
            {8'h00}, /* 0x1c7d */
            {8'h00}, /* 0x1c7c */
            {8'h00}, /* 0x1c7b */
            {8'h00}, /* 0x1c7a */
            {8'h00}, /* 0x1c79 */
            {8'h00}, /* 0x1c78 */
            {8'h00}, /* 0x1c77 */
            {8'h00}, /* 0x1c76 */
            {8'h00}, /* 0x1c75 */
            {8'h00}, /* 0x1c74 */
            {8'h00}, /* 0x1c73 */
            {8'h00}, /* 0x1c72 */
            {8'h00}, /* 0x1c71 */
            {8'h00}, /* 0x1c70 */
            {8'h00}, /* 0x1c6f */
            {8'h00}, /* 0x1c6e */
            {8'h00}, /* 0x1c6d */
            {8'h00}, /* 0x1c6c */
            {8'h00}, /* 0x1c6b */
            {8'h00}, /* 0x1c6a */
            {8'h00}, /* 0x1c69 */
            {8'h00}, /* 0x1c68 */
            {8'h00}, /* 0x1c67 */
            {8'h00}, /* 0x1c66 */
            {8'h00}, /* 0x1c65 */
            {8'h00}, /* 0x1c64 */
            {8'h00}, /* 0x1c63 */
            {8'h00}, /* 0x1c62 */
            {8'h00}, /* 0x1c61 */
            {8'h00}, /* 0x1c60 */
            {8'h00}, /* 0x1c5f */
            {8'h00}, /* 0x1c5e */
            {8'h00}, /* 0x1c5d */
            {8'h00}, /* 0x1c5c */
            {8'h00}, /* 0x1c5b */
            {8'h00}, /* 0x1c5a */
            {8'h00}, /* 0x1c59 */
            {8'h00}, /* 0x1c58 */
            {8'h00}, /* 0x1c57 */
            {8'h00}, /* 0x1c56 */
            {8'h00}, /* 0x1c55 */
            {8'h00}, /* 0x1c54 */
            {8'h00}, /* 0x1c53 */
            {8'h00}, /* 0x1c52 */
            {8'h00}, /* 0x1c51 */
            {8'h00}, /* 0x1c50 */
            {8'h00}, /* 0x1c4f */
            {8'h00}, /* 0x1c4e */
            {8'h00}, /* 0x1c4d */
            {8'h00}, /* 0x1c4c */
            {8'h00}, /* 0x1c4b */
            {8'h00}, /* 0x1c4a */
            {8'h00}, /* 0x1c49 */
            {8'h00}, /* 0x1c48 */
            {8'h00}, /* 0x1c47 */
            {8'h00}, /* 0x1c46 */
            {8'h00}, /* 0x1c45 */
            {8'h00}, /* 0x1c44 */
            {8'h00}, /* 0x1c43 */
            {8'h00}, /* 0x1c42 */
            {8'h00}, /* 0x1c41 */
            {8'h00}, /* 0x1c40 */
            {8'h00}, /* 0x1c3f */
            {8'h00}, /* 0x1c3e */
            {8'h00}, /* 0x1c3d */
            {8'h00}, /* 0x1c3c */
            {8'h00}, /* 0x1c3b */
            {8'h00}, /* 0x1c3a */
            {8'h00}, /* 0x1c39 */
            {8'h00}, /* 0x1c38 */
            {8'h00}, /* 0x1c37 */
            {8'h00}, /* 0x1c36 */
            {8'h00}, /* 0x1c35 */
            {8'h00}, /* 0x1c34 */
            {8'h00}, /* 0x1c33 */
            {8'h00}, /* 0x1c32 */
            {8'h00}, /* 0x1c31 */
            {8'h00}, /* 0x1c30 */
            {8'h00}, /* 0x1c2f */
            {8'h00}, /* 0x1c2e */
            {8'h00}, /* 0x1c2d */
            {8'h00}, /* 0x1c2c */
            {8'h00}, /* 0x1c2b */
            {8'h00}, /* 0x1c2a */
            {8'h00}, /* 0x1c29 */
            {8'h00}, /* 0x1c28 */
            {8'h00}, /* 0x1c27 */
            {8'h00}, /* 0x1c26 */
            {8'h00}, /* 0x1c25 */
            {8'h00}, /* 0x1c24 */
            {8'h00}, /* 0x1c23 */
            {8'h00}, /* 0x1c22 */
            {8'h00}, /* 0x1c21 */
            {8'h00}, /* 0x1c20 */
            {8'h00}, /* 0x1c1f */
            {8'h00}, /* 0x1c1e */
            {8'h00}, /* 0x1c1d */
            {8'h00}, /* 0x1c1c */
            {8'h00}, /* 0x1c1b */
            {8'h00}, /* 0x1c1a */
            {8'h00}, /* 0x1c19 */
            {8'h00}, /* 0x1c18 */
            {8'h00}, /* 0x1c17 */
            {8'h00}, /* 0x1c16 */
            {8'h00}, /* 0x1c15 */
            {8'h00}, /* 0x1c14 */
            {8'h00}, /* 0x1c13 */
            {8'h00}, /* 0x1c12 */
            {8'h00}, /* 0x1c11 */
            {8'h00}, /* 0x1c10 */
            {8'h00}, /* 0x1c0f */
            {8'h00}, /* 0x1c0e */
            {8'h00}, /* 0x1c0d */
            {8'h00}, /* 0x1c0c */
            {8'h00}, /* 0x1c0b */
            {8'h00}, /* 0x1c0a */
            {8'h00}, /* 0x1c09 */
            {8'h00}, /* 0x1c08 */
            {8'h00}, /* 0x1c07 */
            {8'h00}, /* 0x1c06 */
            {8'h00}, /* 0x1c05 */
            {8'h00}, /* 0x1c04 */
            {8'h00}, /* 0x1c03 */
            {8'h00}, /* 0x1c02 */
            {8'h00}, /* 0x1c01 */
            {8'h00}, /* 0x1c00 */
            {8'h00}, /* 0x1bff */
            {8'h00}, /* 0x1bfe */
            {8'h00}, /* 0x1bfd */
            {8'h00}, /* 0x1bfc */
            {8'h00}, /* 0x1bfb */
            {8'h00}, /* 0x1bfa */
            {8'h00}, /* 0x1bf9 */
            {8'h00}, /* 0x1bf8 */
            {8'h00}, /* 0x1bf7 */
            {8'h00}, /* 0x1bf6 */
            {8'h00}, /* 0x1bf5 */
            {8'h00}, /* 0x1bf4 */
            {8'h00}, /* 0x1bf3 */
            {8'h00}, /* 0x1bf2 */
            {8'h00}, /* 0x1bf1 */
            {8'h00}, /* 0x1bf0 */
            {8'h00}, /* 0x1bef */
            {8'h00}, /* 0x1bee */
            {8'h00}, /* 0x1bed */
            {8'h00}, /* 0x1bec */
            {8'h00}, /* 0x1beb */
            {8'h00}, /* 0x1bea */
            {8'h00}, /* 0x1be9 */
            {8'h00}, /* 0x1be8 */
            {8'h00}, /* 0x1be7 */
            {8'h00}, /* 0x1be6 */
            {8'h00}, /* 0x1be5 */
            {8'h00}, /* 0x1be4 */
            {8'h00}, /* 0x1be3 */
            {8'h00}, /* 0x1be2 */
            {8'h00}, /* 0x1be1 */
            {8'h00}, /* 0x1be0 */
            {8'h00}, /* 0x1bdf */
            {8'h00}, /* 0x1bde */
            {8'h00}, /* 0x1bdd */
            {8'h00}, /* 0x1bdc */
            {8'h00}, /* 0x1bdb */
            {8'h00}, /* 0x1bda */
            {8'h00}, /* 0x1bd9 */
            {8'h00}, /* 0x1bd8 */
            {8'h00}, /* 0x1bd7 */
            {8'h00}, /* 0x1bd6 */
            {8'h00}, /* 0x1bd5 */
            {8'h00}, /* 0x1bd4 */
            {8'h00}, /* 0x1bd3 */
            {8'h00}, /* 0x1bd2 */
            {8'h00}, /* 0x1bd1 */
            {8'h00}, /* 0x1bd0 */
            {8'h00}, /* 0x1bcf */
            {8'h00}, /* 0x1bce */
            {8'h00}, /* 0x1bcd */
            {8'h00}, /* 0x1bcc */
            {8'h00}, /* 0x1bcb */
            {8'h00}, /* 0x1bca */
            {8'h00}, /* 0x1bc9 */
            {8'h00}, /* 0x1bc8 */
            {8'h00}, /* 0x1bc7 */
            {8'h00}, /* 0x1bc6 */
            {8'h00}, /* 0x1bc5 */
            {8'h00}, /* 0x1bc4 */
            {8'h00}, /* 0x1bc3 */
            {8'h00}, /* 0x1bc2 */
            {8'h00}, /* 0x1bc1 */
            {8'h00}, /* 0x1bc0 */
            {8'h00}, /* 0x1bbf */
            {8'h00}, /* 0x1bbe */
            {8'h00}, /* 0x1bbd */
            {8'h00}, /* 0x1bbc */
            {8'h00}, /* 0x1bbb */
            {8'h00}, /* 0x1bba */
            {8'h00}, /* 0x1bb9 */
            {8'h00}, /* 0x1bb8 */
            {8'h00}, /* 0x1bb7 */
            {8'h00}, /* 0x1bb6 */
            {8'h00}, /* 0x1bb5 */
            {8'h00}, /* 0x1bb4 */
            {8'h00}, /* 0x1bb3 */
            {8'h00}, /* 0x1bb2 */
            {8'h00}, /* 0x1bb1 */
            {8'h00}, /* 0x1bb0 */
            {8'h00}, /* 0x1baf */
            {8'h00}, /* 0x1bae */
            {8'h00}, /* 0x1bad */
            {8'h00}, /* 0x1bac */
            {8'h00}, /* 0x1bab */
            {8'h00}, /* 0x1baa */
            {8'h00}, /* 0x1ba9 */
            {8'h00}, /* 0x1ba8 */
            {8'h00}, /* 0x1ba7 */
            {8'h00}, /* 0x1ba6 */
            {8'h00}, /* 0x1ba5 */
            {8'h00}, /* 0x1ba4 */
            {8'h00}, /* 0x1ba3 */
            {8'h00}, /* 0x1ba2 */
            {8'h00}, /* 0x1ba1 */
            {8'h00}, /* 0x1ba0 */
            {8'h00}, /* 0x1b9f */
            {8'h00}, /* 0x1b9e */
            {8'h00}, /* 0x1b9d */
            {8'h00}, /* 0x1b9c */
            {8'h00}, /* 0x1b9b */
            {8'h00}, /* 0x1b9a */
            {8'h00}, /* 0x1b99 */
            {8'h00}, /* 0x1b98 */
            {8'h00}, /* 0x1b97 */
            {8'h00}, /* 0x1b96 */
            {8'h00}, /* 0x1b95 */
            {8'h00}, /* 0x1b94 */
            {8'h00}, /* 0x1b93 */
            {8'h00}, /* 0x1b92 */
            {8'h00}, /* 0x1b91 */
            {8'h00}, /* 0x1b90 */
            {8'h00}, /* 0x1b8f */
            {8'h00}, /* 0x1b8e */
            {8'h00}, /* 0x1b8d */
            {8'h00}, /* 0x1b8c */
            {8'h00}, /* 0x1b8b */
            {8'h00}, /* 0x1b8a */
            {8'h00}, /* 0x1b89 */
            {8'h00}, /* 0x1b88 */
            {8'h00}, /* 0x1b87 */
            {8'h00}, /* 0x1b86 */
            {8'h00}, /* 0x1b85 */
            {8'h00}, /* 0x1b84 */
            {8'h00}, /* 0x1b83 */
            {8'h00}, /* 0x1b82 */
            {8'h00}, /* 0x1b81 */
            {8'h00}, /* 0x1b80 */
            {8'h00}, /* 0x1b7f */
            {8'h00}, /* 0x1b7e */
            {8'h00}, /* 0x1b7d */
            {8'h00}, /* 0x1b7c */
            {8'h00}, /* 0x1b7b */
            {8'h00}, /* 0x1b7a */
            {8'h00}, /* 0x1b79 */
            {8'h00}, /* 0x1b78 */
            {8'h00}, /* 0x1b77 */
            {8'h00}, /* 0x1b76 */
            {8'h00}, /* 0x1b75 */
            {8'h00}, /* 0x1b74 */
            {8'h00}, /* 0x1b73 */
            {8'h00}, /* 0x1b72 */
            {8'h00}, /* 0x1b71 */
            {8'h00}, /* 0x1b70 */
            {8'h00}, /* 0x1b6f */
            {8'h00}, /* 0x1b6e */
            {8'h00}, /* 0x1b6d */
            {8'h00}, /* 0x1b6c */
            {8'h00}, /* 0x1b6b */
            {8'h00}, /* 0x1b6a */
            {8'h00}, /* 0x1b69 */
            {8'h00}, /* 0x1b68 */
            {8'h00}, /* 0x1b67 */
            {8'h00}, /* 0x1b66 */
            {8'h00}, /* 0x1b65 */
            {8'h00}, /* 0x1b64 */
            {8'h00}, /* 0x1b63 */
            {8'h00}, /* 0x1b62 */
            {8'h00}, /* 0x1b61 */
            {8'h00}, /* 0x1b60 */
            {8'h00}, /* 0x1b5f */
            {8'h00}, /* 0x1b5e */
            {8'h00}, /* 0x1b5d */
            {8'h00}, /* 0x1b5c */
            {8'h00}, /* 0x1b5b */
            {8'h00}, /* 0x1b5a */
            {8'h00}, /* 0x1b59 */
            {8'h00}, /* 0x1b58 */
            {8'h00}, /* 0x1b57 */
            {8'h00}, /* 0x1b56 */
            {8'h00}, /* 0x1b55 */
            {8'h00}, /* 0x1b54 */
            {8'h00}, /* 0x1b53 */
            {8'h00}, /* 0x1b52 */
            {8'h00}, /* 0x1b51 */
            {8'h00}, /* 0x1b50 */
            {8'h00}, /* 0x1b4f */
            {8'h00}, /* 0x1b4e */
            {8'h00}, /* 0x1b4d */
            {8'h00}, /* 0x1b4c */
            {8'h00}, /* 0x1b4b */
            {8'h00}, /* 0x1b4a */
            {8'h00}, /* 0x1b49 */
            {8'h00}, /* 0x1b48 */
            {8'h00}, /* 0x1b47 */
            {8'h00}, /* 0x1b46 */
            {8'h00}, /* 0x1b45 */
            {8'h00}, /* 0x1b44 */
            {8'h00}, /* 0x1b43 */
            {8'h00}, /* 0x1b42 */
            {8'h00}, /* 0x1b41 */
            {8'h00}, /* 0x1b40 */
            {8'h00}, /* 0x1b3f */
            {8'h00}, /* 0x1b3e */
            {8'h00}, /* 0x1b3d */
            {8'h00}, /* 0x1b3c */
            {8'h00}, /* 0x1b3b */
            {8'h00}, /* 0x1b3a */
            {8'h00}, /* 0x1b39 */
            {8'h00}, /* 0x1b38 */
            {8'h00}, /* 0x1b37 */
            {8'h00}, /* 0x1b36 */
            {8'h00}, /* 0x1b35 */
            {8'h00}, /* 0x1b34 */
            {8'h00}, /* 0x1b33 */
            {8'h00}, /* 0x1b32 */
            {8'h00}, /* 0x1b31 */
            {8'h00}, /* 0x1b30 */
            {8'h00}, /* 0x1b2f */
            {8'h00}, /* 0x1b2e */
            {8'h00}, /* 0x1b2d */
            {8'h00}, /* 0x1b2c */
            {8'h00}, /* 0x1b2b */
            {8'h00}, /* 0x1b2a */
            {8'h00}, /* 0x1b29 */
            {8'h00}, /* 0x1b28 */
            {8'h00}, /* 0x1b27 */
            {8'h00}, /* 0x1b26 */
            {8'h00}, /* 0x1b25 */
            {8'h00}, /* 0x1b24 */
            {8'h00}, /* 0x1b23 */
            {8'h00}, /* 0x1b22 */
            {8'h00}, /* 0x1b21 */
            {8'h00}, /* 0x1b20 */
            {8'h00}, /* 0x1b1f */
            {8'h00}, /* 0x1b1e */
            {8'h00}, /* 0x1b1d */
            {8'h00}, /* 0x1b1c */
            {8'h00}, /* 0x1b1b */
            {8'h00}, /* 0x1b1a */
            {8'h00}, /* 0x1b19 */
            {8'h00}, /* 0x1b18 */
            {8'h00}, /* 0x1b17 */
            {8'h00}, /* 0x1b16 */
            {8'h00}, /* 0x1b15 */
            {8'h00}, /* 0x1b14 */
            {8'h00}, /* 0x1b13 */
            {8'h00}, /* 0x1b12 */
            {8'h00}, /* 0x1b11 */
            {8'h00}, /* 0x1b10 */
            {8'h00}, /* 0x1b0f */
            {8'h00}, /* 0x1b0e */
            {8'h00}, /* 0x1b0d */
            {8'h00}, /* 0x1b0c */
            {8'h00}, /* 0x1b0b */
            {8'h00}, /* 0x1b0a */
            {8'h00}, /* 0x1b09 */
            {8'h00}, /* 0x1b08 */
            {8'h00}, /* 0x1b07 */
            {8'h00}, /* 0x1b06 */
            {8'h00}, /* 0x1b05 */
            {8'h00}, /* 0x1b04 */
            {8'h00}, /* 0x1b03 */
            {8'h00}, /* 0x1b02 */
            {8'h00}, /* 0x1b01 */
            {8'h00}, /* 0x1b00 */
            {8'h00}, /* 0x1aff */
            {8'h00}, /* 0x1afe */
            {8'h00}, /* 0x1afd */
            {8'h00}, /* 0x1afc */
            {8'h00}, /* 0x1afb */
            {8'h00}, /* 0x1afa */
            {8'h00}, /* 0x1af9 */
            {8'h00}, /* 0x1af8 */
            {8'h00}, /* 0x1af7 */
            {8'h00}, /* 0x1af6 */
            {8'h00}, /* 0x1af5 */
            {8'h00}, /* 0x1af4 */
            {8'h00}, /* 0x1af3 */
            {8'h00}, /* 0x1af2 */
            {8'h00}, /* 0x1af1 */
            {8'h00}, /* 0x1af0 */
            {8'h00}, /* 0x1aef */
            {8'h00}, /* 0x1aee */
            {8'h00}, /* 0x1aed */
            {8'h00}, /* 0x1aec */
            {8'h00}, /* 0x1aeb */
            {8'h00}, /* 0x1aea */
            {8'h00}, /* 0x1ae9 */
            {8'h00}, /* 0x1ae8 */
            {8'h00}, /* 0x1ae7 */
            {8'h00}, /* 0x1ae6 */
            {8'h00}, /* 0x1ae5 */
            {8'h00}, /* 0x1ae4 */
            {8'h00}, /* 0x1ae3 */
            {8'h00}, /* 0x1ae2 */
            {8'h00}, /* 0x1ae1 */
            {8'h00}, /* 0x1ae0 */
            {8'h00}, /* 0x1adf */
            {8'h00}, /* 0x1ade */
            {8'h00}, /* 0x1add */
            {8'h00}, /* 0x1adc */
            {8'h00}, /* 0x1adb */
            {8'h00}, /* 0x1ada */
            {8'h00}, /* 0x1ad9 */
            {8'h00}, /* 0x1ad8 */
            {8'h00}, /* 0x1ad7 */
            {8'h00}, /* 0x1ad6 */
            {8'h00}, /* 0x1ad5 */
            {8'h00}, /* 0x1ad4 */
            {8'h00}, /* 0x1ad3 */
            {8'h00}, /* 0x1ad2 */
            {8'h00}, /* 0x1ad1 */
            {8'h00}, /* 0x1ad0 */
            {8'h00}, /* 0x1acf */
            {8'h00}, /* 0x1ace */
            {8'h00}, /* 0x1acd */
            {8'h00}, /* 0x1acc */
            {8'h00}, /* 0x1acb */
            {8'h00}, /* 0x1aca */
            {8'h00}, /* 0x1ac9 */
            {8'h00}, /* 0x1ac8 */
            {8'h00}, /* 0x1ac7 */
            {8'h00}, /* 0x1ac6 */
            {8'h00}, /* 0x1ac5 */
            {8'h00}, /* 0x1ac4 */
            {8'h00}, /* 0x1ac3 */
            {8'h00}, /* 0x1ac2 */
            {8'h00}, /* 0x1ac1 */
            {8'h00}, /* 0x1ac0 */
            {8'h00}, /* 0x1abf */
            {8'h00}, /* 0x1abe */
            {8'h00}, /* 0x1abd */
            {8'h00}, /* 0x1abc */
            {8'h00}, /* 0x1abb */
            {8'h00}, /* 0x1aba */
            {8'h00}, /* 0x1ab9 */
            {8'h00}, /* 0x1ab8 */
            {8'h00}, /* 0x1ab7 */
            {8'h00}, /* 0x1ab6 */
            {8'h00}, /* 0x1ab5 */
            {8'h00}, /* 0x1ab4 */
            {8'h00}, /* 0x1ab3 */
            {8'h00}, /* 0x1ab2 */
            {8'h00}, /* 0x1ab1 */
            {8'h00}, /* 0x1ab0 */
            {8'h00}, /* 0x1aaf */
            {8'h00}, /* 0x1aae */
            {8'h00}, /* 0x1aad */
            {8'h00}, /* 0x1aac */
            {8'h00}, /* 0x1aab */
            {8'h00}, /* 0x1aaa */
            {8'h00}, /* 0x1aa9 */
            {8'h00}, /* 0x1aa8 */
            {8'h00}, /* 0x1aa7 */
            {8'h00}, /* 0x1aa6 */
            {8'h00}, /* 0x1aa5 */
            {8'h00}, /* 0x1aa4 */
            {8'h00}, /* 0x1aa3 */
            {8'h00}, /* 0x1aa2 */
            {8'h00}, /* 0x1aa1 */
            {8'h00}, /* 0x1aa0 */
            {8'h00}, /* 0x1a9f */
            {8'h00}, /* 0x1a9e */
            {8'h00}, /* 0x1a9d */
            {8'h00}, /* 0x1a9c */
            {8'h00}, /* 0x1a9b */
            {8'h00}, /* 0x1a9a */
            {8'h00}, /* 0x1a99 */
            {8'h00}, /* 0x1a98 */
            {8'h00}, /* 0x1a97 */
            {8'h00}, /* 0x1a96 */
            {8'h00}, /* 0x1a95 */
            {8'h00}, /* 0x1a94 */
            {8'h00}, /* 0x1a93 */
            {8'h00}, /* 0x1a92 */
            {8'h00}, /* 0x1a91 */
            {8'h00}, /* 0x1a90 */
            {8'h00}, /* 0x1a8f */
            {8'h00}, /* 0x1a8e */
            {8'h00}, /* 0x1a8d */
            {8'h00}, /* 0x1a8c */
            {8'h00}, /* 0x1a8b */
            {8'h00}, /* 0x1a8a */
            {8'h00}, /* 0x1a89 */
            {8'h00}, /* 0x1a88 */
            {8'h00}, /* 0x1a87 */
            {8'h00}, /* 0x1a86 */
            {8'h00}, /* 0x1a85 */
            {8'h00}, /* 0x1a84 */
            {8'h00}, /* 0x1a83 */
            {8'h00}, /* 0x1a82 */
            {8'h00}, /* 0x1a81 */
            {8'h00}, /* 0x1a80 */
            {8'h00}, /* 0x1a7f */
            {8'h00}, /* 0x1a7e */
            {8'h00}, /* 0x1a7d */
            {8'h00}, /* 0x1a7c */
            {8'h00}, /* 0x1a7b */
            {8'h00}, /* 0x1a7a */
            {8'h00}, /* 0x1a79 */
            {8'h00}, /* 0x1a78 */
            {8'h00}, /* 0x1a77 */
            {8'h00}, /* 0x1a76 */
            {8'h00}, /* 0x1a75 */
            {8'h00}, /* 0x1a74 */
            {8'h00}, /* 0x1a73 */
            {8'h00}, /* 0x1a72 */
            {8'h00}, /* 0x1a71 */
            {8'h00}, /* 0x1a70 */
            {8'h00}, /* 0x1a6f */
            {8'h00}, /* 0x1a6e */
            {8'h00}, /* 0x1a6d */
            {8'h00}, /* 0x1a6c */
            {8'h00}, /* 0x1a6b */
            {8'h00}, /* 0x1a6a */
            {8'h00}, /* 0x1a69 */
            {8'h00}, /* 0x1a68 */
            {8'h00}, /* 0x1a67 */
            {8'h00}, /* 0x1a66 */
            {8'h00}, /* 0x1a65 */
            {8'h00}, /* 0x1a64 */
            {8'h00}, /* 0x1a63 */
            {8'h00}, /* 0x1a62 */
            {8'h00}, /* 0x1a61 */
            {8'h00}, /* 0x1a60 */
            {8'h00}, /* 0x1a5f */
            {8'h00}, /* 0x1a5e */
            {8'h00}, /* 0x1a5d */
            {8'h00}, /* 0x1a5c */
            {8'h00}, /* 0x1a5b */
            {8'h00}, /* 0x1a5a */
            {8'h00}, /* 0x1a59 */
            {8'h00}, /* 0x1a58 */
            {8'h00}, /* 0x1a57 */
            {8'h00}, /* 0x1a56 */
            {8'h00}, /* 0x1a55 */
            {8'h00}, /* 0x1a54 */
            {8'h00}, /* 0x1a53 */
            {8'h00}, /* 0x1a52 */
            {8'h00}, /* 0x1a51 */
            {8'h00}, /* 0x1a50 */
            {8'h00}, /* 0x1a4f */
            {8'h00}, /* 0x1a4e */
            {8'h00}, /* 0x1a4d */
            {8'h00}, /* 0x1a4c */
            {8'h00}, /* 0x1a4b */
            {8'h00}, /* 0x1a4a */
            {8'h00}, /* 0x1a49 */
            {8'h00}, /* 0x1a48 */
            {8'h00}, /* 0x1a47 */
            {8'h00}, /* 0x1a46 */
            {8'h00}, /* 0x1a45 */
            {8'h00}, /* 0x1a44 */
            {8'h00}, /* 0x1a43 */
            {8'h00}, /* 0x1a42 */
            {8'h00}, /* 0x1a41 */
            {8'h00}, /* 0x1a40 */
            {8'h00}, /* 0x1a3f */
            {8'h00}, /* 0x1a3e */
            {8'h00}, /* 0x1a3d */
            {8'h00}, /* 0x1a3c */
            {8'h00}, /* 0x1a3b */
            {8'h00}, /* 0x1a3a */
            {8'h00}, /* 0x1a39 */
            {8'h00}, /* 0x1a38 */
            {8'h00}, /* 0x1a37 */
            {8'h00}, /* 0x1a36 */
            {8'h00}, /* 0x1a35 */
            {8'h00}, /* 0x1a34 */
            {8'h00}, /* 0x1a33 */
            {8'h00}, /* 0x1a32 */
            {8'h00}, /* 0x1a31 */
            {8'h00}, /* 0x1a30 */
            {8'h00}, /* 0x1a2f */
            {8'h00}, /* 0x1a2e */
            {8'h00}, /* 0x1a2d */
            {8'h00}, /* 0x1a2c */
            {8'h00}, /* 0x1a2b */
            {8'h00}, /* 0x1a2a */
            {8'h00}, /* 0x1a29 */
            {8'h00}, /* 0x1a28 */
            {8'h00}, /* 0x1a27 */
            {8'h00}, /* 0x1a26 */
            {8'h00}, /* 0x1a25 */
            {8'h00}, /* 0x1a24 */
            {8'h00}, /* 0x1a23 */
            {8'h00}, /* 0x1a22 */
            {8'h00}, /* 0x1a21 */
            {8'h00}, /* 0x1a20 */
            {8'h00}, /* 0x1a1f */
            {8'h00}, /* 0x1a1e */
            {8'h00}, /* 0x1a1d */
            {8'h00}, /* 0x1a1c */
            {8'h00}, /* 0x1a1b */
            {8'h00}, /* 0x1a1a */
            {8'h00}, /* 0x1a19 */
            {8'h00}, /* 0x1a18 */
            {8'h00}, /* 0x1a17 */
            {8'h00}, /* 0x1a16 */
            {8'h00}, /* 0x1a15 */
            {8'h00}, /* 0x1a14 */
            {8'h00}, /* 0x1a13 */
            {8'h00}, /* 0x1a12 */
            {8'h00}, /* 0x1a11 */
            {8'h00}, /* 0x1a10 */
            {8'h00}, /* 0x1a0f */
            {8'h00}, /* 0x1a0e */
            {8'h00}, /* 0x1a0d */
            {8'h00}, /* 0x1a0c */
            {8'h00}, /* 0x1a0b */
            {8'h00}, /* 0x1a0a */
            {8'h00}, /* 0x1a09 */
            {8'h00}, /* 0x1a08 */
            {8'h00}, /* 0x1a07 */
            {8'h00}, /* 0x1a06 */
            {8'h00}, /* 0x1a05 */
            {8'h00}, /* 0x1a04 */
            {8'h00}, /* 0x1a03 */
            {8'h00}, /* 0x1a02 */
            {8'h00}, /* 0x1a01 */
            {8'h00}, /* 0x1a00 */
            {8'h00}, /* 0x19ff */
            {8'h00}, /* 0x19fe */
            {8'h00}, /* 0x19fd */
            {8'h00}, /* 0x19fc */
            {8'h00}, /* 0x19fb */
            {8'h00}, /* 0x19fa */
            {8'h00}, /* 0x19f9 */
            {8'h00}, /* 0x19f8 */
            {8'h00}, /* 0x19f7 */
            {8'h00}, /* 0x19f6 */
            {8'h00}, /* 0x19f5 */
            {8'h00}, /* 0x19f4 */
            {8'h00}, /* 0x19f3 */
            {8'h00}, /* 0x19f2 */
            {8'h00}, /* 0x19f1 */
            {8'h00}, /* 0x19f0 */
            {8'h00}, /* 0x19ef */
            {8'h00}, /* 0x19ee */
            {8'h00}, /* 0x19ed */
            {8'h00}, /* 0x19ec */
            {8'h00}, /* 0x19eb */
            {8'h00}, /* 0x19ea */
            {8'h00}, /* 0x19e9 */
            {8'h00}, /* 0x19e8 */
            {8'h00}, /* 0x19e7 */
            {8'h00}, /* 0x19e6 */
            {8'h00}, /* 0x19e5 */
            {8'h00}, /* 0x19e4 */
            {8'h00}, /* 0x19e3 */
            {8'h00}, /* 0x19e2 */
            {8'h00}, /* 0x19e1 */
            {8'h00}, /* 0x19e0 */
            {8'h00}, /* 0x19df */
            {8'h00}, /* 0x19de */
            {8'h00}, /* 0x19dd */
            {8'h00}, /* 0x19dc */
            {8'h00}, /* 0x19db */
            {8'h00}, /* 0x19da */
            {8'h00}, /* 0x19d9 */
            {8'h00}, /* 0x19d8 */
            {8'h00}, /* 0x19d7 */
            {8'h00}, /* 0x19d6 */
            {8'h00}, /* 0x19d5 */
            {8'h00}, /* 0x19d4 */
            {8'h00}, /* 0x19d3 */
            {8'h00}, /* 0x19d2 */
            {8'h00}, /* 0x19d1 */
            {8'h00}, /* 0x19d0 */
            {8'h00}, /* 0x19cf */
            {8'h00}, /* 0x19ce */
            {8'h00}, /* 0x19cd */
            {8'h00}, /* 0x19cc */
            {8'h00}, /* 0x19cb */
            {8'h00}, /* 0x19ca */
            {8'h00}, /* 0x19c9 */
            {8'h00}, /* 0x19c8 */
            {8'h00}, /* 0x19c7 */
            {8'h00}, /* 0x19c6 */
            {8'h00}, /* 0x19c5 */
            {8'h00}, /* 0x19c4 */
            {8'h00}, /* 0x19c3 */
            {8'h00}, /* 0x19c2 */
            {8'h00}, /* 0x19c1 */
            {8'h00}, /* 0x19c0 */
            {8'h00}, /* 0x19bf */
            {8'h00}, /* 0x19be */
            {8'h00}, /* 0x19bd */
            {8'h00}, /* 0x19bc */
            {8'h00}, /* 0x19bb */
            {8'h00}, /* 0x19ba */
            {8'h00}, /* 0x19b9 */
            {8'h00}, /* 0x19b8 */
            {8'h00}, /* 0x19b7 */
            {8'h00}, /* 0x19b6 */
            {8'h00}, /* 0x19b5 */
            {8'h00}, /* 0x19b4 */
            {8'h00}, /* 0x19b3 */
            {8'h00}, /* 0x19b2 */
            {8'h00}, /* 0x19b1 */
            {8'h00}, /* 0x19b0 */
            {8'h00}, /* 0x19af */
            {8'h00}, /* 0x19ae */
            {8'h00}, /* 0x19ad */
            {8'h00}, /* 0x19ac */
            {8'h00}, /* 0x19ab */
            {8'h00}, /* 0x19aa */
            {8'h00}, /* 0x19a9 */
            {8'h00}, /* 0x19a8 */
            {8'h00}, /* 0x19a7 */
            {8'h00}, /* 0x19a6 */
            {8'h00}, /* 0x19a5 */
            {8'h00}, /* 0x19a4 */
            {8'h00}, /* 0x19a3 */
            {8'h00}, /* 0x19a2 */
            {8'h00}, /* 0x19a1 */
            {8'h00}, /* 0x19a0 */
            {8'h00}, /* 0x199f */
            {8'h00}, /* 0x199e */
            {8'h00}, /* 0x199d */
            {8'h00}, /* 0x199c */
            {8'h00}, /* 0x199b */
            {8'h00}, /* 0x199a */
            {8'h00}, /* 0x1999 */
            {8'h00}, /* 0x1998 */
            {8'h00}, /* 0x1997 */
            {8'h00}, /* 0x1996 */
            {8'h00}, /* 0x1995 */
            {8'h00}, /* 0x1994 */
            {8'h00}, /* 0x1993 */
            {8'h00}, /* 0x1992 */
            {8'h00}, /* 0x1991 */
            {8'h00}, /* 0x1990 */
            {8'h00}, /* 0x198f */
            {8'h00}, /* 0x198e */
            {8'h00}, /* 0x198d */
            {8'h00}, /* 0x198c */
            {8'h00}, /* 0x198b */
            {8'h00}, /* 0x198a */
            {8'h00}, /* 0x1989 */
            {8'h00}, /* 0x1988 */
            {8'h00}, /* 0x1987 */
            {8'h00}, /* 0x1986 */
            {8'h00}, /* 0x1985 */
            {8'h00}, /* 0x1984 */
            {8'h00}, /* 0x1983 */
            {8'h00}, /* 0x1982 */
            {8'h00}, /* 0x1981 */
            {8'h00}, /* 0x1980 */
            {8'h00}, /* 0x197f */
            {8'h00}, /* 0x197e */
            {8'h00}, /* 0x197d */
            {8'h00}, /* 0x197c */
            {8'h00}, /* 0x197b */
            {8'h00}, /* 0x197a */
            {8'h00}, /* 0x1979 */
            {8'h00}, /* 0x1978 */
            {8'h00}, /* 0x1977 */
            {8'h00}, /* 0x1976 */
            {8'h00}, /* 0x1975 */
            {8'h00}, /* 0x1974 */
            {8'h00}, /* 0x1973 */
            {8'h00}, /* 0x1972 */
            {8'h00}, /* 0x1971 */
            {8'h00}, /* 0x1970 */
            {8'h00}, /* 0x196f */
            {8'h00}, /* 0x196e */
            {8'h00}, /* 0x196d */
            {8'h00}, /* 0x196c */
            {8'h00}, /* 0x196b */
            {8'h00}, /* 0x196a */
            {8'h00}, /* 0x1969 */
            {8'h00}, /* 0x1968 */
            {8'h00}, /* 0x1967 */
            {8'h00}, /* 0x1966 */
            {8'h00}, /* 0x1965 */
            {8'h00}, /* 0x1964 */
            {8'h00}, /* 0x1963 */
            {8'h00}, /* 0x1962 */
            {8'h00}, /* 0x1961 */
            {8'h00}, /* 0x1960 */
            {8'h00}, /* 0x195f */
            {8'h00}, /* 0x195e */
            {8'h00}, /* 0x195d */
            {8'h00}, /* 0x195c */
            {8'h00}, /* 0x195b */
            {8'h00}, /* 0x195a */
            {8'h00}, /* 0x1959 */
            {8'h00}, /* 0x1958 */
            {8'h00}, /* 0x1957 */
            {8'h00}, /* 0x1956 */
            {8'h00}, /* 0x1955 */
            {8'h00}, /* 0x1954 */
            {8'h00}, /* 0x1953 */
            {8'h00}, /* 0x1952 */
            {8'h00}, /* 0x1951 */
            {8'h00}, /* 0x1950 */
            {8'h00}, /* 0x194f */
            {8'h00}, /* 0x194e */
            {8'h00}, /* 0x194d */
            {8'h00}, /* 0x194c */
            {8'h00}, /* 0x194b */
            {8'h00}, /* 0x194a */
            {8'h00}, /* 0x1949 */
            {8'h00}, /* 0x1948 */
            {8'h00}, /* 0x1947 */
            {8'h00}, /* 0x1946 */
            {8'h00}, /* 0x1945 */
            {8'h00}, /* 0x1944 */
            {8'h00}, /* 0x1943 */
            {8'h00}, /* 0x1942 */
            {8'h00}, /* 0x1941 */
            {8'h00}, /* 0x1940 */
            {8'h00}, /* 0x193f */
            {8'h00}, /* 0x193e */
            {8'h00}, /* 0x193d */
            {8'h00}, /* 0x193c */
            {8'h00}, /* 0x193b */
            {8'h00}, /* 0x193a */
            {8'h00}, /* 0x1939 */
            {8'h00}, /* 0x1938 */
            {8'h00}, /* 0x1937 */
            {8'h00}, /* 0x1936 */
            {8'h00}, /* 0x1935 */
            {8'h00}, /* 0x1934 */
            {8'h00}, /* 0x1933 */
            {8'h00}, /* 0x1932 */
            {8'h00}, /* 0x1931 */
            {8'h00}, /* 0x1930 */
            {8'h00}, /* 0x192f */
            {8'h00}, /* 0x192e */
            {8'h00}, /* 0x192d */
            {8'h00}, /* 0x192c */
            {8'h00}, /* 0x192b */
            {8'h00}, /* 0x192a */
            {8'h00}, /* 0x1929 */
            {8'h00}, /* 0x1928 */
            {8'h00}, /* 0x1927 */
            {8'h00}, /* 0x1926 */
            {8'h00}, /* 0x1925 */
            {8'h00}, /* 0x1924 */
            {8'h00}, /* 0x1923 */
            {8'h00}, /* 0x1922 */
            {8'h00}, /* 0x1921 */
            {8'h00}, /* 0x1920 */
            {8'h00}, /* 0x191f */
            {8'h00}, /* 0x191e */
            {8'h00}, /* 0x191d */
            {8'h00}, /* 0x191c */
            {8'h00}, /* 0x191b */
            {8'h00}, /* 0x191a */
            {8'h00}, /* 0x1919 */
            {8'h00}, /* 0x1918 */
            {8'h00}, /* 0x1917 */
            {8'h00}, /* 0x1916 */
            {8'h00}, /* 0x1915 */
            {8'h00}, /* 0x1914 */
            {8'h00}, /* 0x1913 */
            {8'h00}, /* 0x1912 */
            {8'h00}, /* 0x1911 */
            {8'h00}, /* 0x1910 */
            {8'h00}, /* 0x190f */
            {8'h00}, /* 0x190e */
            {8'h00}, /* 0x190d */
            {8'h00}, /* 0x190c */
            {8'h00}, /* 0x190b */
            {8'h00}, /* 0x190a */
            {8'h00}, /* 0x1909 */
            {8'h00}, /* 0x1908 */
            {8'h00}, /* 0x1907 */
            {8'h00}, /* 0x1906 */
            {8'h00}, /* 0x1905 */
            {8'h00}, /* 0x1904 */
            {8'h00}, /* 0x1903 */
            {8'h00}, /* 0x1902 */
            {8'h00}, /* 0x1901 */
            {8'h00}, /* 0x1900 */
            {8'h00}, /* 0x18ff */
            {8'h00}, /* 0x18fe */
            {8'h00}, /* 0x18fd */
            {8'h00}, /* 0x18fc */
            {8'h00}, /* 0x18fb */
            {8'h00}, /* 0x18fa */
            {8'h00}, /* 0x18f9 */
            {8'h00}, /* 0x18f8 */
            {8'h00}, /* 0x18f7 */
            {8'h00}, /* 0x18f6 */
            {8'h00}, /* 0x18f5 */
            {8'h00}, /* 0x18f4 */
            {8'h00}, /* 0x18f3 */
            {8'h00}, /* 0x18f2 */
            {8'h00}, /* 0x18f1 */
            {8'h00}, /* 0x18f0 */
            {8'h00}, /* 0x18ef */
            {8'h00}, /* 0x18ee */
            {8'h00}, /* 0x18ed */
            {8'h00}, /* 0x18ec */
            {8'h00}, /* 0x18eb */
            {8'h00}, /* 0x18ea */
            {8'h00}, /* 0x18e9 */
            {8'h00}, /* 0x18e8 */
            {8'h00}, /* 0x18e7 */
            {8'h00}, /* 0x18e6 */
            {8'h00}, /* 0x18e5 */
            {8'h00}, /* 0x18e4 */
            {8'h00}, /* 0x18e3 */
            {8'h00}, /* 0x18e2 */
            {8'h00}, /* 0x18e1 */
            {8'h00}, /* 0x18e0 */
            {8'h00}, /* 0x18df */
            {8'h00}, /* 0x18de */
            {8'h00}, /* 0x18dd */
            {8'h00}, /* 0x18dc */
            {8'h00}, /* 0x18db */
            {8'h00}, /* 0x18da */
            {8'h00}, /* 0x18d9 */
            {8'h00}, /* 0x18d8 */
            {8'h00}, /* 0x18d7 */
            {8'h00}, /* 0x18d6 */
            {8'h00}, /* 0x18d5 */
            {8'h00}, /* 0x18d4 */
            {8'h00}, /* 0x18d3 */
            {8'h00}, /* 0x18d2 */
            {8'h00}, /* 0x18d1 */
            {8'h00}, /* 0x18d0 */
            {8'h00}, /* 0x18cf */
            {8'h00}, /* 0x18ce */
            {8'h00}, /* 0x18cd */
            {8'h00}, /* 0x18cc */
            {8'h00}, /* 0x18cb */
            {8'h00}, /* 0x18ca */
            {8'h00}, /* 0x18c9 */
            {8'h00}, /* 0x18c8 */
            {8'h00}, /* 0x18c7 */
            {8'h00}, /* 0x18c6 */
            {8'h00}, /* 0x18c5 */
            {8'h00}, /* 0x18c4 */
            {8'h00}, /* 0x18c3 */
            {8'h00}, /* 0x18c2 */
            {8'h00}, /* 0x18c1 */
            {8'h00}, /* 0x18c0 */
            {8'h00}, /* 0x18bf */
            {8'h00}, /* 0x18be */
            {8'h00}, /* 0x18bd */
            {8'h00}, /* 0x18bc */
            {8'h00}, /* 0x18bb */
            {8'h00}, /* 0x18ba */
            {8'h00}, /* 0x18b9 */
            {8'h00}, /* 0x18b8 */
            {8'h00}, /* 0x18b7 */
            {8'h00}, /* 0x18b6 */
            {8'h00}, /* 0x18b5 */
            {8'h00}, /* 0x18b4 */
            {8'h00}, /* 0x18b3 */
            {8'h00}, /* 0x18b2 */
            {8'h00}, /* 0x18b1 */
            {8'h00}, /* 0x18b0 */
            {8'h00}, /* 0x18af */
            {8'h00}, /* 0x18ae */
            {8'h00}, /* 0x18ad */
            {8'h00}, /* 0x18ac */
            {8'h00}, /* 0x18ab */
            {8'h00}, /* 0x18aa */
            {8'h00}, /* 0x18a9 */
            {8'h00}, /* 0x18a8 */
            {8'h00}, /* 0x18a7 */
            {8'h00}, /* 0x18a6 */
            {8'h00}, /* 0x18a5 */
            {8'h00}, /* 0x18a4 */
            {8'h00}, /* 0x18a3 */
            {8'h00}, /* 0x18a2 */
            {8'h00}, /* 0x18a1 */
            {8'h00}, /* 0x18a0 */
            {8'h00}, /* 0x189f */
            {8'h00}, /* 0x189e */
            {8'h00}, /* 0x189d */
            {8'h00}, /* 0x189c */
            {8'h00}, /* 0x189b */
            {8'h00}, /* 0x189a */
            {8'h00}, /* 0x1899 */
            {8'h00}, /* 0x1898 */
            {8'h00}, /* 0x1897 */
            {8'h00}, /* 0x1896 */
            {8'h00}, /* 0x1895 */
            {8'h00}, /* 0x1894 */
            {8'h00}, /* 0x1893 */
            {8'h00}, /* 0x1892 */
            {8'h00}, /* 0x1891 */
            {8'h00}, /* 0x1890 */
            {8'h00}, /* 0x188f */
            {8'h00}, /* 0x188e */
            {8'h00}, /* 0x188d */
            {8'h00}, /* 0x188c */
            {8'h00}, /* 0x188b */
            {8'h00}, /* 0x188a */
            {8'h00}, /* 0x1889 */
            {8'h00}, /* 0x1888 */
            {8'h00}, /* 0x1887 */
            {8'h00}, /* 0x1886 */
            {8'h00}, /* 0x1885 */
            {8'h00}, /* 0x1884 */
            {8'h00}, /* 0x1883 */
            {8'h00}, /* 0x1882 */
            {8'h00}, /* 0x1881 */
            {8'h00}, /* 0x1880 */
            {8'h00}, /* 0x187f */
            {8'h00}, /* 0x187e */
            {8'h00}, /* 0x187d */
            {8'h00}, /* 0x187c */
            {8'h00}, /* 0x187b */
            {8'h00}, /* 0x187a */
            {8'h00}, /* 0x1879 */
            {8'h00}, /* 0x1878 */
            {8'h00}, /* 0x1877 */
            {8'h00}, /* 0x1876 */
            {8'h00}, /* 0x1875 */
            {8'h00}, /* 0x1874 */
            {8'h00}, /* 0x1873 */
            {8'h00}, /* 0x1872 */
            {8'h00}, /* 0x1871 */
            {8'h00}, /* 0x1870 */
            {8'h00}, /* 0x186f */
            {8'h00}, /* 0x186e */
            {8'h00}, /* 0x186d */
            {8'h00}, /* 0x186c */
            {8'h00}, /* 0x186b */
            {8'h00}, /* 0x186a */
            {8'h00}, /* 0x1869 */
            {8'h00}, /* 0x1868 */
            {8'h00}, /* 0x1867 */
            {8'h00}, /* 0x1866 */
            {8'h00}, /* 0x1865 */
            {8'h00}, /* 0x1864 */
            {8'h00}, /* 0x1863 */
            {8'h00}, /* 0x1862 */
            {8'h00}, /* 0x1861 */
            {8'h00}, /* 0x1860 */
            {8'h00}, /* 0x185f */
            {8'h00}, /* 0x185e */
            {8'h00}, /* 0x185d */
            {8'h00}, /* 0x185c */
            {8'h00}, /* 0x185b */
            {8'h00}, /* 0x185a */
            {8'h00}, /* 0x1859 */
            {8'h00}, /* 0x1858 */
            {8'h00}, /* 0x1857 */
            {8'h00}, /* 0x1856 */
            {8'h00}, /* 0x1855 */
            {8'h00}, /* 0x1854 */
            {8'h00}, /* 0x1853 */
            {8'h00}, /* 0x1852 */
            {8'h00}, /* 0x1851 */
            {8'h00}, /* 0x1850 */
            {8'h00}, /* 0x184f */
            {8'h00}, /* 0x184e */
            {8'h00}, /* 0x184d */
            {8'h00}, /* 0x184c */
            {8'h00}, /* 0x184b */
            {8'h00}, /* 0x184a */
            {8'h00}, /* 0x1849 */
            {8'h00}, /* 0x1848 */
            {8'h00}, /* 0x1847 */
            {8'h00}, /* 0x1846 */
            {8'h00}, /* 0x1845 */
            {8'h00}, /* 0x1844 */
            {8'h00}, /* 0x1843 */
            {8'h00}, /* 0x1842 */
            {8'h00}, /* 0x1841 */
            {8'h00}, /* 0x1840 */
            {8'h00}, /* 0x183f */
            {8'h00}, /* 0x183e */
            {8'h00}, /* 0x183d */
            {8'h00}, /* 0x183c */
            {8'h00}, /* 0x183b */
            {8'h00}, /* 0x183a */
            {8'h00}, /* 0x1839 */
            {8'h00}, /* 0x1838 */
            {8'h00}, /* 0x1837 */
            {8'h00}, /* 0x1836 */
            {8'h00}, /* 0x1835 */
            {8'h00}, /* 0x1834 */
            {8'h00}, /* 0x1833 */
            {8'h00}, /* 0x1832 */
            {8'h00}, /* 0x1831 */
            {8'h00}, /* 0x1830 */
            {8'h00}, /* 0x182f */
            {8'h00}, /* 0x182e */
            {8'h00}, /* 0x182d */
            {8'h00}, /* 0x182c */
            {8'h00}, /* 0x182b */
            {8'h00}, /* 0x182a */
            {8'h00}, /* 0x1829 */
            {8'h00}, /* 0x1828 */
            {8'h00}, /* 0x1827 */
            {8'h00}, /* 0x1826 */
            {8'h00}, /* 0x1825 */
            {8'h00}, /* 0x1824 */
            {8'h00}, /* 0x1823 */
            {8'h00}, /* 0x1822 */
            {8'h00}, /* 0x1821 */
            {8'h00}, /* 0x1820 */
            {8'h00}, /* 0x181f */
            {8'h00}, /* 0x181e */
            {8'h00}, /* 0x181d */
            {8'h00}, /* 0x181c */
            {8'h00}, /* 0x181b */
            {8'h00}, /* 0x181a */
            {8'h00}, /* 0x1819 */
            {8'h00}, /* 0x1818 */
            {8'h00}, /* 0x1817 */
            {8'h00}, /* 0x1816 */
            {8'h00}, /* 0x1815 */
            {8'h00}, /* 0x1814 */
            {8'h00}, /* 0x1813 */
            {8'h00}, /* 0x1812 */
            {8'h00}, /* 0x1811 */
            {8'h00}, /* 0x1810 */
            {8'h00}, /* 0x180f */
            {8'h00}, /* 0x180e */
            {8'h00}, /* 0x180d */
            {8'h00}, /* 0x180c */
            {8'h00}, /* 0x180b */
            {8'h00}, /* 0x180a */
            {8'h00}, /* 0x1809 */
            {8'h00}, /* 0x1808 */
            {8'h00}, /* 0x1807 */
            {8'h00}, /* 0x1806 */
            {8'h00}, /* 0x1805 */
            {8'h00}, /* 0x1804 */
            {8'h00}, /* 0x1803 */
            {8'h00}, /* 0x1802 */
            {8'h00}, /* 0x1801 */
            {8'h00}, /* 0x1800 */
            {8'h00}, /* 0x17ff */
            {8'h00}, /* 0x17fe */
            {8'h00}, /* 0x17fd */
            {8'h00}, /* 0x17fc */
            {8'h00}, /* 0x17fb */
            {8'h00}, /* 0x17fa */
            {8'h00}, /* 0x17f9 */
            {8'h00}, /* 0x17f8 */
            {8'h00}, /* 0x17f7 */
            {8'h00}, /* 0x17f6 */
            {8'h00}, /* 0x17f5 */
            {8'h00}, /* 0x17f4 */
            {8'h00}, /* 0x17f3 */
            {8'h00}, /* 0x17f2 */
            {8'h00}, /* 0x17f1 */
            {8'h00}, /* 0x17f0 */
            {8'h00}, /* 0x17ef */
            {8'h00}, /* 0x17ee */
            {8'h00}, /* 0x17ed */
            {8'h00}, /* 0x17ec */
            {8'h00}, /* 0x17eb */
            {8'h00}, /* 0x17ea */
            {8'h00}, /* 0x17e9 */
            {8'h00}, /* 0x17e8 */
            {8'h00}, /* 0x17e7 */
            {8'h00}, /* 0x17e6 */
            {8'h00}, /* 0x17e5 */
            {8'h00}, /* 0x17e4 */
            {8'h00}, /* 0x17e3 */
            {8'h00}, /* 0x17e2 */
            {8'h00}, /* 0x17e1 */
            {8'h00}, /* 0x17e0 */
            {8'h00}, /* 0x17df */
            {8'h00}, /* 0x17de */
            {8'h00}, /* 0x17dd */
            {8'h00}, /* 0x17dc */
            {8'h00}, /* 0x17db */
            {8'h00}, /* 0x17da */
            {8'h00}, /* 0x17d9 */
            {8'h00}, /* 0x17d8 */
            {8'h00}, /* 0x17d7 */
            {8'h00}, /* 0x17d6 */
            {8'h00}, /* 0x17d5 */
            {8'h00}, /* 0x17d4 */
            {8'h00}, /* 0x17d3 */
            {8'h00}, /* 0x17d2 */
            {8'h00}, /* 0x17d1 */
            {8'h00}, /* 0x17d0 */
            {8'h00}, /* 0x17cf */
            {8'h00}, /* 0x17ce */
            {8'h00}, /* 0x17cd */
            {8'h00}, /* 0x17cc */
            {8'h00}, /* 0x17cb */
            {8'h00}, /* 0x17ca */
            {8'h00}, /* 0x17c9 */
            {8'h00}, /* 0x17c8 */
            {8'h00}, /* 0x17c7 */
            {8'h00}, /* 0x17c6 */
            {8'h00}, /* 0x17c5 */
            {8'h00}, /* 0x17c4 */
            {8'h00}, /* 0x17c3 */
            {8'h00}, /* 0x17c2 */
            {8'h00}, /* 0x17c1 */
            {8'h00}, /* 0x17c0 */
            {8'h00}, /* 0x17bf */
            {8'h00}, /* 0x17be */
            {8'h00}, /* 0x17bd */
            {8'h00}, /* 0x17bc */
            {8'h00}, /* 0x17bb */
            {8'h00}, /* 0x17ba */
            {8'h00}, /* 0x17b9 */
            {8'h00}, /* 0x17b8 */
            {8'h00}, /* 0x17b7 */
            {8'h00}, /* 0x17b6 */
            {8'h00}, /* 0x17b5 */
            {8'h00}, /* 0x17b4 */
            {8'h00}, /* 0x17b3 */
            {8'h00}, /* 0x17b2 */
            {8'h00}, /* 0x17b1 */
            {8'h00}, /* 0x17b0 */
            {8'h00}, /* 0x17af */
            {8'h00}, /* 0x17ae */
            {8'h00}, /* 0x17ad */
            {8'h00}, /* 0x17ac */
            {8'h00}, /* 0x17ab */
            {8'h00}, /* 0x17aa */
            {8'h00}, /* 0x17a9 */
            {8'h00}, /* 0x17a8 */
            {8'h00}, /* 0x17a7 */
            {8'h00}, /* 0x17a6 */
            {8'h00}, /* 0x17a5 */
            {8'h00}, /* 0x17a4 */
            {8'h00}, /* 0x17a3 */
            {8'h00}, /* 0x17a2 */
            {8'h00}, /* 0x17a1 */
            {8'h00}, /* 0x17a0 */
            {8'h00}, /* 0x179f */
            {8'h00}, /* 0x179e */
            {8'h00}, /* 0x179d */
            {8'h00}, /* 0x179c */
            {8'h00}, /* 0x179b */
            {8'h00}, /* 0x179a */
            {8'h00}, /* 0x1799 */
            {8'h00}, /* 0x1798 */
            {8'h00}, /* 0x1797 */
            {8'h00}, /* 0x1796 */
            {8'h00}, /* 0x1795 */
            {8'h00}, /* 0x1794 */
            {8'h00}, /* 0x1793 */
            {8'h00}, /* 0x1792 */
            {8'h00}, /* 0x1791 */
            {8'h00}, /* 0x1790 */
            {8'h00}, /* 0x178f */
            {8'h00}, /* 0x178e */
            {8'h00}, /* 0x178d */
            {8'h00}, /* 0x178c */
            {8'h00}, /* 0x178b */
            {8'h00}, /* 0x178a */
            {8'h00}, /* 0x1789 */
            {8'h00}, /* 0x1788 */
            {8'h00}, /* 0x1787 */
            {8'h00}, /* 0x1786 */
            {8'h00}, /* 0x1785 */
            {8'h00}, /* 0x1784 */
            {8'h00}, /* 0x1783 */
            {8'h00}, /* 0x1782 */
            {8'h00}, /* 0x1781 */
            {8'h00}, /* 0x1780 */
            {8'h00}, /* 0x177f */
            {8'h00}, /* 0x177e */
            {8'h00}, /* 0x177d */
            {8'h00}, /* 0x177c */
            {8'h00}, /* 0x177b */
            {8'h00}, /* 0x177a */
            {8'h00}, /* 0x1779 */
            {8'h00}, /* 0x1778 */
            {8'h00}, /* 0x1777 */
            {8'h00}, /* 0x1776 */
            {8'h00}, /* 0x1775 */
            {8'h00}, /* 0x1774 */
            {8'h00}, /* 0x1773 */
            {8'h00}, /* 0x1772 */
            {8'h00}, /* 0x1771 */
            {8'h00}, /* 0x1770 */
            {8'h00}, /* 0x176f */
            {8'h00}, /* 0x176e */
            {8'h00}, /* 0x176d */
            {8'h00}, /* 0x176c */
            {8'h00}, /* 0x176b */
            {8'h00}, /* 0x176a */
            {8'h00}, /* 0x1769 */
            {8'h00}, /* 0x1768 */
            {8'h00}, /* 0x1767 */
            {8'h00}, /* 0x1766 */
            {8'h00}, /* 0x1765 */
            {8'h00}, /* 0x1764 */
            {8'h00}, /* 0x1763 */
            {8'h00}, /* 0x1762 */
            {8'h00}, /* 0x1761 */
            {8'h00}, /* 0x1760 */
            {8'h00}, /* 0x175f */
            {8'h00}, /* 0x175e */
            {8'h00}, /* 0x175d */
            {8'h00}, /* 0x175c */
            {8'h00}, /* 0x175b */
            {8'h00}, /* 0x175a */
            {8'h00}, /* 0x1759 */
            {8'h00}, /* 0x1758 */
            {8'h00}, /* 0x1757 */
            {8'h00}, /* 0x1756 */
            {8'h00}, /* 0x1755 */
            {8'h00}, /* 0x1754 */
            {8'h00}, /* 0x1753 */
            {8'h00}, /* 0x1752 */
            {8'h00}, /* 0x1751 */
            {8'h00}, /* 0x1750 */
            {8'h00}, /* 0x174f */
            {8'h00}, /* 0x174e */
            {8'h00}, /* 0x174d */
            {8'h00}, /* 0x174c */
            {8'h00}, /* 0x174b */
            {8'h00}, /* 0x174a */
            {8'h00}, /* 0x1749 */
            {8'h00}, /* 0x1748 */
            {8'h00}, /* 0x1747 */
            {8'h00}, /* 0x1746 */
            {8'h00}, /* 0x1745 */
            {8'h00}, /* 0x1744 */
            {8'h00}, /* 0x1743 */
            {8'h00}, /* 0x1742 */
            {8'h00}, /* 0x1741 */
            {8'h00}, /* 0x1740 */
            {8'h00}, /* 0x173f */
            {8'h00}, /* 0x173e */
            {8'h00}, /* 0x173d */
            {8'h00}, /* 0x173c */
            {8'h00}, /* 0x173b */
            {8'h00}, /* 0x173a */
            {8'h00}, /* 0x1739 */
            {8'h00}, /* 0x1738 */
            {8'h00}, /* 0x1737 */
            {8'h00}, /* 0x1736 */
            {8'h00}, /* 0x1735 */
            {8'h00}, /* 0x1734 */
            {8'h00}, /* 0x1733 */
            {8'h00}, /* 0x1732 */
            {8'h00}, /* 0x1731 */
            {8'h00}, /* 0x1730 */
            {8'h00}, /* 0x172f */
            {8'h00}, /* 0x172e */
            {8'h00}, /* 0x172d */
            {8'h00}, /* 0x172c */
            {8'h00}, /* 0x172b */
            {8'h00}, /* 0x172a */
            {8'h00}, /* 0x1729 */
            {8'h00}, /* 0x1728 */
            {8'h00}, /* 0x1727 */
            {8'h00}, /* 0x1726 */
            {8'h00}, /* 0x1725 */
            {8'h00}, /* 0x1724 */
            {8'h00}, /* 0x1723 */
            {8'h00}, /* 0x1722 */
            {8'h00}, /* 0x1721 */
            {8'h00}, /* 0x1720 */
            {8'h00}, /* 0x171f */
            {8'h00}, /* 0x171e */
            {8'h00}, /* 0x171d */
            {8'h00}, /* 0x171c */
            {8'h00}, /* 0x171b */
            {8'h00}, /* 0x171a */
            {8'h00}, /* 0x1719 */
            {8'h00}, /* 0x1718 */
            {8'h00}, /* 0x1717 */
            {8'h00}, /* 0x1716 */
            {8'h00}, /* 0x1715 */
            {8'h00}, /* 0x1714 */
            {8'h00}, /* 0x1713 */
            {8'h00}, /* 0x1712 */
            {8'h00}, /* 0x1711 */
            {8'h00}, /* 0x1710 */
            {8'h00}, /* 0x170f */
            {8'h00}, /* 0x170e */
            {8'h00}, /* 0x170d */
            {8'h00}, /* 0x170c */
            {8'h00}, /* 0x170b */
            {8'h00}, /* 0x170a */
            {8'h00}, /* 0x1709 */
            {8'h00}, /* 0x1708 */
            {8'h00}, /* 0x1707 */
            {8'h00}, /* 0x1706 */
            {8'h00}, /* 0x1705 */
            {8'h00}, /* 0x1704 */
            {8'h00}, /* 0x1703 */
            {8'h00}, /* 0x1702 */
            {8'h00}, /* 0x1701 */
            {8'h00}, /* 0x1700 */
            {8'h00}, /* 0x16ff */
            {8'h00}, /* 0x16fe */
            {8'h00}, /* 0x16fd */
            {8'h00}, /* 0x16fc */
            {8'h00}, /* 0x16fb */
            {8'h00}, /* 0x16fa */
            {8'h00}, /* 0x16f9 */
            {8'h00}, /* 0x16f8 */
            {8'h00}, /* 0x16f7 */
            {8'h00}, /* 0x16f6 */
            {8'h00}, /* 0x16f5 */
            {8'h00}, /* 0x16f4 */
            {8'h00}, /* 0x16f3 */
            {8'h00}, /* 0x16f2 */
            {8'h00}, /* 0x16f1 */
            {8'h00}, /* 0x16f0 */
            {8'h00}, /* 0x16ef */
            {8'h00}, /* 0x16ee */
            {8'h00}, /* 0x16ed */
            {8'h00}, /* 0x16ec */
            {8'h00}, /* 0x16eb */
            {8'h00}, /* 0x16ea */
            {8'h00}, /* 0x16e9 */
            {8'h00}, /* 0x16e8 */
            {8'h00}, /* 0x16e7 */
            {8'h00}, /* 0x16e6 */
            {8'h00}, /* 0x16e5 */
            {8'h00}, /* 0x16e4 */
            {8'h00}, /* 0x16e3 */
            {8'h00}, /* 0x16e2 */
            {8'h00}, /* 0x16e1 */
            {8'h00}, /* 0x16e0 */
            {8'h00}, /* 0x16df */
            {8'h00}, /* 0x16de */
            {8'h00}, /* 0x16dd */
            {8'h00}, /* 0x16dc */
            {8'h00}, /* 0x16db */
            {8'h00}, /* 0x16da */
            {8'h00}, /* 0x16d9 */
            {8'h00}, /* 0x16d8 */
            {8'h00}, /* 0x16d7 */
            {8'h00}, /* 0x16d6 */
            {8'h00}, /* 0x16d5 */
            {8'h00}, /* 0x16d4 */
            {8'h00}, /* 0x16d3 */
            {8'h00}, /* 0x16d2 */
            {8'h00}, /* 0x16d1 */
            {8'h00}, /* 0x16d0 */
            {8'h00}, /* 0x16cf */
            {8'h00}, /* 0x16ce */
            {8'h00}, /* 0x16cd */
            {8'h00}, /* 0x16cc */
            {8'h00}, /* 0x16cb */
            {8'h00}, /* 0x16ca */
            {8'h00}, /* 0x16c9 */
            {8'h00}, /* 0x16c8 */
            {8'h00}, /* 0x16c7 */
            {8'h00}, /* 0x16c6 */
            {8'h00}, /* 0x16c5 */
            {8'h00}, /* 0x16c4 */
            {8'h00}, /* 0x16c3 */
            {8'h00}, /* 0x16c2 */
            {8'h00}, /* 0x16c1 */
            {8'h00}, /* 0x16c0 */
            {8'h00}, /* 0x16bf */
            {8'h00}, /* 0x16be */
            {8'h00}, /* 0x16bd */
            {8'h00}, /* 0x16bc */
            {8'h00}, /* 0x16bb */
            {8'h00}, /* 0x16ba */
            {8'h00}, /* 0x16b9 */
            {8'h00}, /* 0x16b8 */
            {8'h00}, /* 0x16b7 */
            {8'h00}, /* 0x16b6 */
            {8'h00}, /* 0x16b5 */
            {8'h00}, /* 0x16b4 */
            {8'h00}, /* 0x16b3 */
            {8'h00}, /* 0x16b2 */
            {8'h00}, /* 0x16b1 */
            {8'h00}, /* 0x16b0 */
            {8'h00}, /* 0x16af */
            {8'h00}, /* 0x16ae */
            {8'h00}, /* 0x16ad */
            {8'h00}, /* 0x16ac */
            {8'h00}, /* 0x16ab */
            {8'h00}, /* 0x16aa */
            {8'h00}, /* 0x16a9 */
            {8'h00}, /* 0x16a8 */
            {8'h00}, /* 0x16a7 */
            {8'h00}, /* 0x16a6 */
            {8'h00}, /* 0x16a5 */
            {8'h00}, /* 0x16a4 */
            {8'h00}, /* 0x16a3 */
            {8'h00}, /* 0x16a2 */
            {8'h00}, /* 0x16a1 */
            {8'h00}, /* 0x16a0 */
            {8'h00}, /* 0x169f */
            {8'h00}, /* 0x169e */
            {8'h00}, /* 0x169d */
            {8'h00}, /* 0x169c */
            {8'h00}, /* 0x169b */
            {8'h00}, /* 0x169a */
            {8'h00}, /* 0x1699 */
            {8'h00}, /* 0x1698 */
            {8'h00}, /* 0x1697 */
            {8'h00}, /* 0x1696 */
            {8'h00}, /* 0x1695 */
            {8'h00}, /* 0x1694 */
            {8'h00}, /* 0x1693 */
            {8'h00}, /* 0x1692 */
            {8'h00}, /* 0x1691 */
            {8'h00}, /* 0x1690 */
            {8'h00}, /* 0x168f */
            {8'h00}, /* 0x168e */
            {8'h00}, /* 0x168d */
            {8'h00}, /* 0x168c */
            {8'h00}, /* 0x168b */
            {8'h00}, /* 0x168a */
            {8'h00}, /* 0x1689 */
            {8'h00}, /* 0x1688 */
            {8'h00}, /* 0x1687 */
            {8'h00}, /* 0x1686 */
            {8'h00}, /* 0x1685 */
            {8'h00}, /* 0x1684 */
            {8'h00}, /* 0x1683 */
            {8'h00}, /* 0x1682 */
            {8'h00}, /* 0x1681 */
            {8'h00}, /* 0x1680 */
            {8'h00}, /* 0x167f */
            {8'h00}, /* 0x167e */
            {8'h00}, /* 0x167d */
            {8'h00}, /* 0x167c */
            {8'h00}, /* 0x167b */
            {8'h00}, /* 0x167a */
            {8'h00}, /* 0x1679 */
            {8'h00}, /* 0x1678 */
            {8'h00}, /* 0x1677 */
            {8'h00}, /* 0x1676 */
            {8'h00}, /* 0x1675 */
            {8'h00}, /* 0x1674 */
            {8'h00}, /* 0x1673 */
            {8'h00}, /* 0x1672 */
            {8'h00}, /* 0x1671 */
            {8'h00}, /* 0x1670 */
            {8'h00}, /* 0x166f */
            {8'h00}, /* 0x166e */
            {8'h00}, /* 0x166d */
            {8'h00}, /* 0x166c */
            {8'h00}, /* 0x166b */
            {8'h00}, /* 0x166a */
            {8'h00}, /* 0x1669 */
            {8'h00}, /* 0x1668 */
            {8'h00}, /* 0x1667 */
            {8'h00}, /* 0x1666 */
            {8'h00}, /* 0x1665 */
            {8'h00}, /* 0x1664 */
            {8'h00}, /* 0x1663 */
            {8'h00}, /* 0x1662 */
            {8'h00}, /* 0x1661 */
            {8'h00}, /* 0x1660 */
            {8'h00}, /* 0x165f */
            {8'h00}, /* 0x165e */
            {8'h00}, /* 0x165d */
            {8'h00}, /* 0x165c */
            {8'h00}, /* 0x165b */
            {8'h00}, /* 0x165a */
            {8'h00}, /* 0x1659 */
            {8'h00}, /* 0x1658 */
            {8'h00}, /* 0x1657 */
            {8'h00}, /* 0x1656 */
            {8'h00}, /* 0x1655 */
            {8'h00}, /* 0x1654 */
            {8'h00}, /* 0x1653 */
            {8'h00}, /* 0x1652 */
            {8'h00}, /* 0x1651 */
            {8'h00}, /* 0x1650 */
            {8'h00}, /* 0x164f */
            {8'h00}, /* 0x164e */
            {8'h00}, /* 0x164d */
            {8'h00}, /* 0x164c */
            {8'h00}, /* 0x164b */
            {8'h00}, /* 0x164a */
            {8'h00}, /* 0x1649 */
            {8'h00}, /* 0x1648 */
            {8'h00}, /* 0x1647 */
            {8'h00}, /* 0x1646 */
            {8'h00}, /* 0x1645 */
            {8'h00}, /* 0x1644 */
            {8'h00}, /* 0x1643 */
            {8'h00}, /* 0x1642 */
            {8'h00}, /* 0x1641 */
            {8'h00}, /* 0x1640 */
            {8'h00}, /* 0x163f */
            {8'h00}, /* 0x163e */
            {8'h00}, /* 0x163d */
            {8'h00}, /* 0x163c */
            {8'h00}, /* 0x163b */
            {8'h00}, /* 0x163a */
            {8'h00}, /* 0x1639 */
            {8'h00}, /* 0x1638 */
            {8'h00}, /* 0x1637 */
            {8'h00}, /* 0x1636 */
            {8'h00}, /* 0x1635 */
            {8'h00}, /* 0x1634 */
            {8'h00}, /* 0x1633 */
            {8'h00}, /* 0x1632 */
            {8'h00}, /* 0x1631 */
            {8'h00}, /* 0x1630 */
            {8'h00}, /* 0x162f */
            {8'h00}, /* 0x162e */
            {8'h00}, /* 0x162d */
            {8'h00}, /* 0x162c */
            {8'h00}, /* 0x162b */
            {8'h00}, /* 0x162a */
            {8'h00}, /* 0x1629 */
            {8'h00}, /* 0x1628 */
            {8'h00}, /* 0x1627 */
            {8'h00}, /* 0x1626 */
            {8'h00}, /* 0x1625 */
            {8'h00}, /* 0x1624 */
            {8'h00}, /* 0x1623 */
            {8'h00}, /* 0x1622 */
            {8'h00}, /* 0x1621 */
            {8'h00}, /* 0x1620 */
            {8'h00}, /* 0x161f */
            {8'h00}, /* 0x161e */
            {8'h00}, /* 0x161d */
            {8'h00}, /* 0x161c */
            {8'h00}, /* 0x161b */
            {8'h00}, /* 0x161a */
            {8'h00}, /* 0x1619 */
            {8'h00}, /* 0x1618 */
            {8'h00}, /* 0x1617 */
            {8'h00}, /* 0x1616 */
            {8'h00}, /* 0x1615 */
            {8'h00}, /* 0x1614 */
            {8'h00}, /* 0x1613 */
            {8'h00}, /* 0x1612 */
            {8'h00}, /* 0x1611 */
            {8'h00}, /* 0x1610 */
            {8'h00}, /* 0x160f */
            {8'h00}, /* 0x160e */
            {8'h00}, /* 0x160d */
            {8'h00}, /* 0x160c */
            {8'h00}, /* 0x160b */
            {8'h00}, /* 0x160a */
            {8'h00}, /* 0x1609 */
            {8'h00}, /* 0x1608 */
            {8'h00}, /* 0x1607 */
            {8'h00}, /* 0x1606 */
            {8'h00}, /* 0x1605 */
            {8'h00}, /* 0x1604 */
            {8'h00}, /* 0x1603 */
            {8'h00}, /* 0x1602 */
            {8'h00}, /* 0x1601 */
            {8'h00}, /* 0x1600 */
            {8'h00}, /* 0x15ff */
            {8'h00}, /* 0x15fe */
            {8'h00}, /* 0x15fd */
            {8'h00}, /* 0x15fc */
            {8'h00}, /* 0x15fb */
            {8'h00}, /* 0x15fa */
            {8'h00}, /* 0x15f9 */
            {8'h00}, /* 0x15f8 */
            {8'h00}, /* 0x15f7 */
            {8'h00}, /* 0x15f6 */
            {8'h00}, /* 0x15f5 */
            {8'h00}, /* 0x15f4 */
            {8'h00}, /* 0x15f3 */
            {8'h00}, /* 0x15f2 */
            {8'h00}, /* 0x15f1 */
            {8'h00}, /* 0x15f0 */
            {8'h00}, /* 0x15ef */
            {8'h00}, /* 0x15ee */
            {8'h00}, /* 0x15ed */
            {8'h00}, /* 0x15ec */
            {8'h00}, /* 0x15eb */
            {8'h00}, /* 0x15ea */
            {8'h00}, /* 0x15e9 */
            {8'h00}, /* 0x15e8 */
            {8'h00}, /* 0x15e7 */
            {8'h00}, /* 0x15e6 */
            {8'h00}, /* 0x15e5 */
            {8'h00}, /* 0x15e4 */
            {8'h00}, /* 0x15e3 */
            {8'h00}, /* 0x15e2 */
            {8'h00}, /* 0x15e1 */
            {8'h00}, /* 0x15e0 */
            {8'h00}, /* 0x15df */
            {8'h00}, /* 0x15de */
            {8'h00}, /* 0x15dd */
            {8'h00}, /* 0x15dc */
            {8'h00}, /* 0x15db */
            {8'h00}, /* 0x15da */
            {8'h00}, /* 0x15d9 */
            {8'h00}, /* 0x15d8 */
            {8'h00}, /* 0x15d7 */
            {8'h00}, /* 0x15d6 */
            {8'h00}, /* 0x15d5 */
            {8'h00}, /* 0x15d4 */
            {8'h00}, /* 0x15d3 */
            {8'h00}, /* 0x15d2 */
            {8'h00}, /* 0x15d1 */
            {8'h00}, /* 0x15d0 */
            {8'h00}, /* 0x15cf */
            {8'h00}, /* 0x15ce */
            {8'h00}, /* 0x15cd */
            {8'h00}, /* 0x15cc */
            {8'h00}, /* 0x15cb */
            {8'h00}, /* 0x15ca */
            {8'h00}, /* 0x15c9 */
            {8'h00}, /* 0x15c8 */
            {8'h00}, /* 0x15c7 */
            {8'h00}, /* 0x15c6 */
            {8'h00}, /* 0x15c5 */
            {8'h00}, /* 0x15c4 */
            {8'h00}, /* 0x15c3 */
            {8'h00}, /* 0x15c2 */
            {8'h00}, /* 0x15c1 */
            {8'h00}, /* 0x15c0 */
            {8'h00}, /* 0x15bf */
            {8'h00}, /* 0x15be */
            {8'h00}, /* 0x15bd */
            {8'h00}, /* 0x15bc */
            {8'h00}, /* 0x15bb */
            {8'h00}, /* 0x15ba */
            {8'h00}, /* 0x15b9 */
            {8'h00}, /* 0x15b8 */
            {8'h00}, /* 0x15b7 */
            {8'h00}, /* 0x15b6 */
            {8'h00}, /* 0x15b5 */
            {8'h00}, /* 0x15b4 */
            {8'h00}, /* 0x15b3 */
            {8'h00}, /* 0x15b2 */
            {8'h00}, /* 0x15b1 */
            {8'h00}, /* 0x15b0 */
            {8'h00}, /* 0x15af */
            {8'h00}, /* 0x15ae */
            {8'h00}, /* 0x15ad */
            {8'h00}, /* 0x15ac */
            {8'h00}, /* 0x15ab */
            {8'h00}, /* 0x15aa */
            {8'h00}, /* 0x15a9 */
            {8'h00}, /* 0x15a8 */
            {8'h00}, /* 0x15a7 */
            {8'h00}, /* 0x15a6 */
            {8'h00}, /* 0x15a5 */
            {8'h00}, /* 0x15a4 */
            {8'h00}, /* 0x15a3 */
            {8'h00}, /* 0x15a2 */
            {8'h00}, /* 0x15a1 */
            {8'h00}, /* 0x15a0 */
            {8'h00}, /* 0x159f */
            {8'h00}, /* 0x159e */
            {8'h00}, /* 0x159d */
            {8'h00}, /* 0x159c */
            {8'h00}, /* 0x159b */
            {8'h00}, /* 0x159a */
            {8'h00}, /* 0x1599 */
            {8'h00}, /* 0x1598 */
            {8'h00}, /* 0x1597 */
            {8'h00}, /* 0x1596 */
            {8'h00}, /* 0x1595 */
            {8'h00}, /* 0x1594 */
            {8'h00}, /* 0x1593 */
            {8'h00}, /* 0x1592 */
            {8'h00}, /* 0x1591 */
            {8'h00}, /* 0x1590 */
            {8'h00}, /* 0x158f */
            {8'h00}, /* 0x158e */
            {8'h00}, /* 0x158d */
            {8'h00}, /* 0x158c */
            {8'h00}, /* 0x158b */
            {8'h00}, /* 0x158a */
            {8'h00}, /* 0x1589 */
            {8'h00}, /* 0x1588 */
            {8'h00}, /* 0x1587 */
            {8'h00}, /* 0x1586 */
            {8'h00}, /* 0x1585 */
            {8'h00}, /* 0x1584 */
            {8'h00}, /* 0x1583 */
            {8'h00}, /* 0x1582 */
            {8'h00}, /* 0x1581 */
            {8'h00}, /* 0x1580 */
            {8'h00}, /* 0x157f */
            {8'h00}, /* 0x157e */
            {8'h00}, /* 0x157d */
            {8'h00}, /* 0x157c */
            {8'h00}, /* 0x157b */
            {8'h00}, /* 0x157a */
            {8'h00}, /* 0x1579 */
            {8'h00}, /* 0x1578 */
            {8'h00}, /* 0x1577 */
            {8'h00}, /* 0x1576 */
            {8'h00}, /* 0x1575 */
            {8'h00}, /* 0x1574 */
            {8'h00}, /* 0x1573 */
            {8'h00}, /* 0x1572 */
            {8'h00}, /* 0x1571 */
            {8'h00}, /* 0x1570 */
            {8'h00}, /* 0x156f */
            {8'h00}, /* 0x156e */
            {8'h00}, /* 0x156d */
            {8'h00}, /* 0x156c */
            {8'h00}, /* 0x156b */
            {8'h00}, /* 0x156a */
            {8'h00}, /* 0x1569 */
            {8'h00}, /* 0x1568 */
            {8'h00}, /* 0x1567 */
            {8'h00}, /* 0x1566 */
            {8'h00}, /* 0x1565 */
            {8'h00}, /* 0x1564 */
            {8'h00}, /* 0x1563 */
            {8'h00}, /* 0x1562 */
            {8'h00}, /* 0x1561 */
            {8'h00}, /* 0x1560 */
            {8'h00}, /* 0x155f */
            {8'h00}, /* 0x155e */
            {8'h00}, /* 0x155d */
            {8'h00}, /* 0x155c */
            {8'h00}, /* 0x155b */
            {8'h00}, /* 0x155a */
            {8'h00}, /* 0x1559 */
            {8'h00}, /* 0x1558 */
            {8'h00}, /* 0x1557 */
            {8'h00}, /* 0x1556 */
            {8'h00}, /* 0x1555 */
            {8'h00}, /* 0x1554 */
            {8'h00}, /* 0x1553 */
            {8'h00}, /* 0x1552 */
            {8'h00}, /* 0x1551 */
            {8'h00}, /* 0x1550 */
            {8'h00}, /* 0x154f */
            {8'h00}, /* 0x154e */
            {8'h00}, /* 0x154d */
            {8'h00}, /* 0x154c */
            {8'h00}, /* 0x154b */
            {8'h00}, /* 0x154a */
            {8'h00}, /* 0x1549 */
            {8'h00}, /* 0x1548 */
            {8'h00}, /* 0x1547 */
            {8'h00}, /* 0x1546 */
            {8'h00}, /* 0x1545 */
            {8'h00}, /* 0x1544 */
            {8'h00}, /* 0x1543 */
            {8'h00}, /* 0x1542 */
            {8'h00}, /* 0x1541 */
            {8'h00}, /* 0x1540 */
            {8'h00}, /* 0x153f */
            {8'h00}, /* 0x153e */
            {8'h00}, /* 0x153d */
            {8'h00}, /* 0x153c */
            {8'h00}, /* 0x153b */
            {8'h00}, /* 0x153a */
            {8'h00}, /* 0x1539 */
            {8'h00}, /* 0x1538 */
            {8'h00}, /* 0x1537 */
            {8'h00}, /* 0x1536 */
            {8'h00}, /* 0x1535 */
            {8'h00}, /* 0x1534 */
            {8'h00}, /* 0x1533 */
            {8'h00}, /* 0x1532 */
            {8'h00}, /* 0x1531 */
            {8'h00}, /* 0x1530 */
            {8'h00}, /* 0x152f */
            {8'h00}, /* 0x152e */
            {8'h00}, /* 0x152d */
            {8'h00}, /* 0x152c */
            {8'h00}, /* 0x152b */
            {8'h00}, /* 0x152a */
            {8'h00}, /* 0x1529 */
            {8'h00}, /* 0x1528 */
            {8'h00}, /* 0x1527 */
            {8'h00}, /* 0x1526 */
            {8'h00}, /* 0x1525 */
            {8'h00}, /* 0x1524 */
            {8'h00}, /* 0x1523 */
            {8'h00}, /* 0x1522 */
            {8'h00}, /* 0x1521 */
            {8'h00}, /* 0x1520 */
            {8'h00}, /* 0x151f */
            {8'h00}, /* 0x151e */
            {8'h00}, /* 0x151d */
            {8'h00}, /* 0x151c */
            {8'h00}, /* 0x151b */
            {8'h00}, /* 0x151a */
            {8'h00}, /* 0x1519 */
            {8'h00}, /* 0x1518 */
            {8'h00}, /* 0x1517 */
            {8'h00}, /* 0x1516 */
            {8'h00}, /* 0x1515 */
            {8'h00}, /* 0x1514 */
            {8'h00}, /* 0x1513 */
            {8'h00}, /* 0x1512 */
            {8'h00}, /* 0x1511 */
            {8'h00}, /* 0x1510 */
            {8'h00}, /* 0x150f */
            {8'h00}, /* 0x150e */
            {8'h00}, /* 0x150d */
            {8'h00}, /* 0x150c */
            {8'h00}, /* 0x150b */
            {8'h00}, /* 0x150a */
            {8'h00}, /* 0x1509 */
            {8'h00}, /* 0x1508 */
            {8'h00}, /* 0x1507 */
            {8'h00}, /* 0x1506 */
            {8'h00}, /* 0x1505 */
            {8'h00}, /* 0x1504 */
            {8'h00}, /* 0x1503 */
            {8'h00}, /* 0x1502 */
            {8'h00}, /* 0x1501 */
            {8'h00}, /* 0x1500 */
            {8'h00}, /* 0x14ff */
            {8'h00}, /* 0x14fe */
            {8'h00}, /* 0x14fd */
            {8'h00}, /* 0x14fc */
            {8'h00}, /* 0x14fb */
            {8'h00}, /* 0x14fa */
            {8'h00}, /* 0x14f9 */
            {8'h00}, /* 0x14f8 */
            {8'h00}, /* 0x14f7 */
            {8'h00}, /* 0x14f6 */
            {8'h00}, /* 0x14f5 */
            {8'h00}, /* 0x14f4 */
            {8'h00}, /* 0x14f3 */
            {8'h00}, /* 0x14f2 */
            {8'h00}, /* 0x14f1 */
            {8'h00}, /* 0x14f0 */
            {8'h00}, /* 0x14ef */
            {8'h00}, /* 0x14ee */
            {8'h00}, /* 0x14ed */
            {8'h00}, /* 0x14ec */
            {8'h00}, /* 0x14eb */
            {8'h00}, /* 0x14ea */
            {8'h00}, /* 0x14e9 */
            {8'h00}, /* 0x14e8 */
            {8'h00}, /* 0x14e7 */
            {8'h00}, /* 0x14e6 */
            {8'h00}, /* 0x14e5 */
            {8'h00}, /* 0x14e4 */
            {8'h00}, /* 0x14e3 */
            {8'h00}, /* 0x14e2 */
            {8'h00}, /* 0x14e1 */
            {8'h00}, /* 0x14e0 */
            {8'h00}, /* 0x14df */
            {8'h00}, /* 0x14de */
            {8'h00}, /* 0x14dd */
            {8'h00}, /* 0x14dc */
            {8'h00}, /* 0x14db */
            {8'h00}, /* 0x14da */
            {8'h00}, /* 0x14d9 */
            {8'h00}, /* 0x14d8 */
            {8'h00}, /* 0x14d7 */
            {8'h00}, /* 0x14d6 */
            {8'h00}, /* 0x14d5 */
            {8'h00}, /* 0x14d4 */
            {8'h00}, /* 0x14d3 */
            {8'h00}, /* 0x14d2 */
            {8'h00}, /* 0x14d1 */
            {8'h00}, /* 0x14d0 */
            {8'h00}, /* 0x14cf */
            {8'h00}, /* 0x14ce */
            {8'h00}, /* 0x14cd */
            {8'h00}, /* 0x14cc */
            {8'h00}, /* 0x14cb */
            {8'h00}, /* 0x14ca */
            {8'h00}, /* 0x14c9 */
            {8'h00}, /* 0x14c8 */
            {8'h00}, /* 0x14c7 */
            {8'h00}, /* 0x14c6 */
            {8'h00}, /* 0x14c5 */
            {8'h00}, /* 0x14c4 */
            {8'h00}, /* 0x14c3 */
            {8'h00}, /* 0x14c2 */
            {8'h00}, /* 0x14c1 */
            {8'h00}, /* 0x14c0 */
            {8'h00}, /* 0x14bf */
            {8'h00}, /* 0x14be */
            {8'h00}, /* 0x14bd */
            {8'h00}, /* 0x14bc */
            {8'h00}, /* 0x14bb */
            {8'h00}, /* 0x14ba */
            {8'h00}, /* 0x14b9 */
            {8'h00}, /* 0x14b8 */
            {8'h00}, /* 0x14b7 */
            {8'h00}, /* 0x14b6 */
            {8'h00}, /* 0x14b5 */
            {8'h00}, /* 0x14b4 */
            {8'h00}, /* 0x14b3 */
            {8'h00}, /* 0x14b2 */
            {8'h00}, /* 0x14b1 */
            {8'h00}, /* 0x14b0 */
            {8'h00}, /* 0x14af */
            {8'h00}, /* 0x14ae */
            {8'h00}, /* 0x14ad */
            {8'h00}, /* 0x14ac */
            {8'h00}, /* 0x14ab */
            {8'h00}, /* 0x14aa */
            {8'h00}, /* 0x14a9 */
            {8'h00}, /* 0x14a8 */
            {8'h00}, /* 0x14a7 */
            {8'h00}, /* 0x14a6 */
            {8'h00}, /* 0x14a5 */
            {8'h00}, /* 0x14a4 */
            {8'h00}, /* 0x14a3 */
            {8'h00}, /* 0x14a2 */
            {8'h00}, /* 0x14a1 */
            {8'h00}, /* 0x14a0 */
            {8'h00}, /* 0x149f */
            {8'h00}, /* 0x149e */
            {8'h00}, /* 0x149d */
            {8'h00}, /* 0x149c */
            {8'h00}, /* 0x149b */
            {8'h00}, /* 0x149a */
            {8'h00}, /* 0x1499 */
            {8'h00}, /* 0x1498 */
            {8'h00}, /* 0x1497 */
            {8'h00}, /* 0x1496 */
            {8'h00}, /* 0x1495 */
            {8'h00}, /* 0x1494 */
            {8'h00}, /* 0x1493 */
            {8'h00}, /* 0x1492 */
            {8'h00}, /* 0x1491 */
            {8'h00}, /* 0x1490 */
            {8'h00}, /* 0x148f */
            {8'h00}, /* 0x148e */
            {8'h00}, /* 0x148d */
            {8'h00}, /* 0x148c */
            {8'h00}, /* 0x148b */
            {8'h00}, /* 0x148a */
            {8'h00}, /* 0x1489 */
            {8'h00}, /* 0x1488 */
            {8'h00}, /* 0x1487 */
            {8'h00}, /* 0x1486 */
            {8'h00}, /* 0x1485 */
            {8'h00}, /* 0x1484 */
            {8'h00}, /* 0x1483 */
            {8'h00}, /* 0x1482 */
            {8'h00}, /* 0x1481 */
            {8'h00}, /* 0x1480 */
            {8'h00}, /* 0x147f */
            {8'h00}, /* 0x147e */
            {8'h00}, /* 0x147d */
            {8'h00}, /* 0x147c */
            {8'h00}, /* 0x147b */
            {8'h00}, /* 0x147a */
            {8'h00}, /* 0x1479 */
            {8'h00}, /* 0x1478 */
            {8'h00}, /* 0x1477 */
            {8'h00}, /* 0x1476 */
            {8'h00}, /* 0x1475 */
            {8'h00}, /* 0x1474 */
            {8'h00}, /* 0x1473 */
            {8'h00}, /* 0x1472 */
            {8'h00}, /* 0x1471 */
            {8'h00}, /* 0x1470 */
            {8'h00}, /* 0x146f */
            {8'h00}, /* 0x146e */
            {8'h00}, /* 0x146d */
            {8'h00}, /* 0x146c */
            {8'h00}, /* 0x146b */
            {8'h00}, /* 0x146a */
            {8'h00}, /* 0x1469 */
            {8'h00}, /* 0x1468 */
            {8'h00}, /* 0x1467 */
            {8'h00}, /* 0x1466 */
            {8'h00}, /* 0x1465 */
            {8'h00}, /* 0x1464 */
            {8'h00}, /* 0x1463 */
            {8'h00}, /* 0x1462 */
            {8'h00}, /* 0x1461 */
            {8'h00}, /* 0x1460 */
            {8'h00}, /* 0x145f */
            {8'h00}, /* 0x145e */
            {8'h00}, /* 0x145d */
            {8'h00}, /* 0x145c */
            {8'h00}, /* 0x145b */
            {8'h00}, /* 0x145a */
            {8'h00}, /* 0x1459 */
            {8'h00}, /* 0x1458 */
            {8'h00}, /* 0x1457 */
            {8'h00}, /* 0x1456 */
            {8'h00}, /* 0x1455 */
            {8'h00}, /* 0x1454 */
            {8'h00}, /* 0x1453 */
            {8'h00}, /* 0x1452 */
            {8'h00}, /* 0x1451 */
            {8'h00}, /* 0x1450 */
            {8'h00}, /* 0x144f */
            {8'h00}, /* 0x144e */
            {8'h00}, /* 0x144d */
            {8'h00}, /* 0x144c */
            {8'h00}, /* 0x144b */
            {8'h00}, /* 0x144a */
            {8'h00}, /* 0x1449 */
            {8'h00}, /* 0x1448 */
            {8'h00}, /* 0x1447 */
            {8'h00}, /* 0x1446 */
            {8'h00}, /* 0x1445 */
            {8'h00}, /* 0x1444 */
            {8'h00}, /* 0x1443 */
            {8'h00}, /* 0x1442 */
            {8'h00}, /* 0x1441 */
            {8'h00}, /* 0x1440 */
            {8'h00}, /* 0x143f */
            {8'h00}, /* 0x143e */
            {8'h00}, /* 0x143d */
            {8'h00}, /* 0x143c */
            {8'h00}, /* 0x143b */
            {8'h00}, /* 0x143a */
            {8'h00}, /* 0x1439 */
            {8'h00}, /* 0x1438 */
            {8'h00}, /* 0x1437 */
            {8'h00}, /* 0x1436 */
            {8'h00}, /* 0x1435 */
            {8'h00}, /* 0x1434 */
            {8'h00}, /* 0x1433 */
            {8'h00}, /* 0x1432 */
            {8'h00}, /* 0x1431 */
            {8'h00}, /* 0x1430 */
            {8'h00}, /* 0x142f */
            {8'h00}, /* 0x142e */
            {8'h00}, /* 0x142d */
            {8'h00}, /* 0x142c */
            {8'h00}, /* 0x142b */
            {8'h00}, /* 0x142a */
            {8'h00}, /* 0x1429 */
            {8'h00}, /* 0x1428 */
            {8'h00}, /* 0x1427 */
            {8'h00}, /* 0x1426 */
            {8'h00}, /* 0x1425 */
            {8'h00}, /* 0x1424 */
            {8'h00}, /* 0x1423 */
            {8'h00}, /* 0x1422 */
            {8'h00}, /* 0x1421 */
            {8'h00}, /* 0x1420 */
            {8'h00}, /* 0x141f */
            {8'h00}, /* 0x141e */
            {8'h00}, /* 0x141d */
            {8'h00}, /* 0x141c */
            {8'h00}, /* 0x141b */
            {8'h00}, /* 0x141a */
            {8'h00}, /* 0x1419 */
            {8'h00}, /* 0x1418 */
            {8'h00}, /* 0x1417 */
            {8'h00}, /* 0x1416 */
            {8'h00}, /* 0x1415 */
            {8'h00}, /* 0x1414 */
            {8'h00}, /* 0x1413 */
            {8'h00}, /* 0x1412 */
            {8'h00}, /* 0x1411 */
            {8'h00}, /* 0x1410 */
            {8'h00}, /* 0x140f */
            {8'h00}, /* 0x140e */
            {8'h00}, /* 0x140d */
            {8'h00}, /* 0x140c */
            {8'h00}, /* 0x140b */
            {8'h00}, /* 0x140a */
            {8'h00}, /* 0x1409 */
            {8'h00}, /* 0x1408 */
            {8'h00}, /* 0x1407 */
            {8'h00}, /* 0x1406 */
            {8'h00}, /* 0x1405 */
            {8'h00}, /* 0x1404 */
            {8'h00}, /* 0x1403 */
            {8'h00}, /* 0x1402 */
            {8'h00}, /* 0x1401 */
            {8'h00}, /* 0x1400 */
            {8'h00}, /* 0x13ff */
            {8'h00}, /* 0x13fe */
            {8'h00}, /* 0x13fd */
            {8'h00}, /* 0x13fc */
            {8'h00}, /* 0x13fb */
            {8'h00}, /* 0x13fa */
            {8'h00}, /* 0x13f9 */
            {8'h00}, /* 0x13f8 */
            {8'h00}, /* 0x13f7 */
            {8'h00}, /* 0x13f6 */
            {8'h00}, /* 0x13f5 */
            {8'h00}, /* 0x13f4 */
            {8'h00}, /* 0x13f3 */
            {8'h00}, /* 0x13f2 */
            {8'h00}, /* 0x13f1 */
            {8'h00}, /* 0x13f0 */
            {8'h00}, /* 0x13ef */
            {8'h00}, /* 0x13ee */
            {8'h00}, /* 0x13ed */
            {8'h00}, /* 0x13ec */
            {8'h00}, /* 0x13eb */
            {8'h00}, /* 0x13ea */
            {8'h00}, /* 0x13e9 */
            {8'h00}, /* 0x13e8 */
            {8'h00}, /* 0x13e7 */
            {8'h00}, /* 0x13e6 */
            {8'h00}, /* 0x13e5 */
            {8'h00}, /* 0x13e4 */
            {8'h00}, /* 0x13e3 */
            {8'h00}, /* 0x13e2 */
            {8'h00}, /* 0x13e1 */
            {8'h00}, /* 0x13e0 */
            {8'h00}, /* 0x13df */
            {8'h00}, /* 0x13de */
            {8'h00}, /* 0x13dd */
            {8'h00}, /* 0x13dc */
            {8'h00}, /* 0x13db */
            {8'h00}, /* 0x13da */
            {8'h00}, /* 0x13d9 */
            {8'h00}, /* 0x13d8 */
            {8'h00}, /* 0x13d7 */
            {8'h00}, /* 0x13d6 */
            {8'h00}, /* 0x13d5 */
            {8'h00}, /* 0x13d4 */
            {8'h00}, /* 0x13d3 */
            {8'h00}, /* 0x13d2 */
            {8'h00}, /* 0x13d1 */
            {8'h00}, /* 0x13d0 */
            {8'h00}, /* 0x13cf */
            {8'h00}, /* 0x13ce */
            {8'h00}, /* 0x13cd */
            {8'h00}, /* 0x13cc */
            {8'h00}, /* 0x13cb */
            {8'h00}, /* 0x13ca */
            {8'h00}, /* 0x13c9 */
            {8'h00}, /* 0x13c8 */
            {8'h00}, /* 0x13c7 */
            {8'h00}, /* 0x13c6 */
            {8'h00}, /* 0x13c5 */
            {8'h00}, /* 0x13c4 */
            {8'h00}, /* 0x13c3 */
            {8'h00}, /* 0x13c2 */
            {8'h00}, /* 0x13c1 */
            {8'h00}, /* 0x13c0 */
            {8'h00}, /* 0x13bf */
            {8'h00}, /* 0x13be */
            {8'h00}, /* 0x13bd */
            {8'h00}, /* 0x13bc */
            {8'h00}, /* 0x13bb */
            {8'h00}, /* 0x13ba */
            {8'h00}, /* 0x13b9 */
            {8'h00}, /* 0x13b8 */
            {8'h00}, /* 0x13b7 */
            {8'h00}, /* 0x13b6 */
            {8'h00}, /* 0x13b5 */
            {8'h00}, /* 0x13b4 */
            {8'h00}, /* 0x13b3 */
            {8'h00}, /* 0x13b2 */
            {8'h00}, /* 0x13b1 */
            {8'h00}, /* 0x13b0 */
            {8'h00}, /* 0x13af */
            {8'h00}, /* 0x13ae */
            {8'h00}, /* 0x13ad */
            {8'h00}, /* 0x13ac */
            {8'h00}, /* 0x13ab */
            {8'h00}, /* 0x13aa */
            {8'h00}, /* 0x13a9 */
            {8'h00}, /* 0x13a8 */
            {8'h00}, /* 0x13a7 */
            {8'h00}, /* 0x13a6 */
            {8'h00}, /* 0x13a5 */
            {8'h00}, /* 0x13a4 */
            {8'h00}, /* 0x13a3 */
            {8'h00}, /* 0x13a2 */
            {8'h00}, /* 0x13a1 */
            {8'h00}, /* 0x13a0 */
            {8'h00}, /* 0x139f */
            {8'h00}, /* 0x139e */
            {8'h00}, /* 0x139d */
            {8'h00}, /* 0x139c */
            {8'h00}, /* 0x139b */
            {8'h00}, /* 0x139a */
            {8'h00}, /* 0x1399 */
            {8'h00}, /* 0x1398 */
            {8'h00}, /* 0x1397 */
            {8'h00}, /* 0x1396 */
            {8'h00}, /* 0x1395 */
            {8'h00}, /* 0x1394 */
            {8'h00}, /* 0x1393 */
            {8'h00}, /* 0x1392 */
            {8'h00}, /* 0x1391 */
            {8'h00}, /* 0x1390 */
            {8'h00}, /* 0x138f */
            {8'h00}, /* 0x138e */
            {8'h00}, /* 0x138d */
            {8'h00}, /* 0x138c */
            {8'h00}, /* 0x138b */
            {8'h00}, /* 0x138a */
            {8'h00}, /* 0x1389 */
            {8'h00}, /* 0x1388 */
            {8'h00}, /* 0x1387 */
            {8'h00}, /* 0x1386 */
            {8'h00}, /* 0x1385 */
            {8'h00}, /* 0x1384 */
            {8'h00}, /* 0x1383 */
            {8'h00}, /* 0x1382 */
            {8'h00}, /* 0x1381 */
            {8'h00}, /* 0x1380 */
            {8'h00}, /* 0x137f */
            {8'h00}, /* 0x137e */
            {8'h00}, /* 0x137d */
            {8'h00}, /* 0x137c */
            {8'h00}, /* 0x137b */
            {8'h00}, /* 0x137a */
            {8'h00}, /* 0x1379 */
            {8'h00}, /* 0x1378 */
            {8'h00}, /* 0x1377 */
            {8'h00}, /* 0x1376 */
            {8'h00}, /* 0x1375 */
            {8'h00}, /* 0x1374 */
            {8'h00}, /* 0x1373 */
            {8'h00}, /* 0x1372 */
            {8'h00}, /* 0x1371 */
            {8'h00}, /* 0x1370 */
            {8'h00}, /* 0x136f */
            {8'h00}, /* 0x136e */
            {8'h00}, /* 0x136d */
            {8'h00}, /* 0x136c */
            {8'h00}, /* 0x136b */
            {8'h00}, /* 0x136a */
            {8'h00}, /* 0x1369 */
            {8'h00}, /* 0x1368 */
            {8'h00}, /* 0x1367 */
            {8'h00}, /* 0x1366 */
            {8'h00}, /* 0x1365 */
            {8'h00}, /* 0x1364 */
            {8'h00}, /* 0x1363 */
            {8'h00}, /* 0x1362 */
            {8'h00}, /* 0x1361 */
            {8'h00}, /* 0x1360 */
            {8'h00}, /* 0x135f */
            {8'h00}, /* 0x135e */
            {8'h00}, /* 0x135d */
            {8'h00}, /* 0x135c */
            {8'h00}, /* 0x135b */
            {8'h00}, /* 0x135a */
            {8'h00}, /* 0x1359 */
            {8'h00}, /* 0x1358 */
            {8'h00}, /* 0x1357 */
            {8'h00}, /* 0x1356 */
            {8'h00}, /* 0x1355 */
            {8'h00}, /* 0x1354 */
            {8'h00}, /* 0x1353 */
            {8'h00}, /* 0x1352 */
            {8'h00}, /* 0x1351 */
            {8'h00}, /* 0x1350 */
            {8'h00}, /* 0x134f */
            {8'h00}, /* 0x134e */
            {8'h00}, /* 0x134d */
            {8'h00}, /* 0x134c */
            {8'h00}, /* 0x134b */
            {8'h00}, /* 0x134a */
            {8'h00}, /* 0x1349 */
            {8'h00}, /* 0x1348 */
            {8'h00}, /* 0x1347 */
            {8'h00}, /* 0x1346 */
            {8'h00}, /* 0x1345 */
            {8'h00}, /* 0x1344 */
            {8'h00}, /* 0x1343 */
            {8'h00}, /* 0x1342 */
            {8'h00}, /* 0x1341 */
            {8'h00}, /* 0x1340 */
            {8'h00}, /* 0x133f */
            {8'h00}, /* 0x133e */
            {8'h00}, /* 0x133d */
            {8'h00}, /* 0x133c */
            {8'h00}, /* 0x133b */
            {8'h00}, /* 0x133a */
            {8'h00}, /* 0x1339 */
            {8'h00}, /* 0x1338 */
            {8'h00}, /* 0x1337 */
            {8'h00}, /* 0x1336 */
            {8'h00}, /* 0x1335 */
            {8'h00}, /* 0x1334 */
            {8'h00}, /* 0x1333 */
            {8'h00}, /* 0x1332 */
            {8'h00}, /* 0x1331 */
            {8'h00}, /* 0x1330 */
            {8'h00}, /* 0x132f */
            {8'h00}, /* 0x132e */
            {8'h00}, /* 0x132d */
            {8'h00}, /* 0x132c */
            {8'h00}, /* 0x132b */
            {8'h00}, /* 0x132a */
            {8'h00}, /* 0x1329 */
            {8'h00}, /* 0x1328 */
            {8'h00}, /* 0x1327 */
            {8'h00}, /* 0x1326 */
            {8'h00}, /* 0x1325 */
            {8'h00}, /* 0x1324 */
            {8'h00}, /* 0x1323 */
            {8'h00}, /* 0x1322 */
            {8'h00}, /* 0x1321 */
            {8'h00}, /* 0x1320 */
            {8'h00}, /* 0x131f */
            {8'h00}, /* 0x131e */
            {8'h00}, /* 0x131d */
            {8'h00}, /* 0x131c */
            {8'h00}, /* 0x131b */
            {8'h00}, /* 0x131a */
            {8'h00}, /* 0x1319 */
            {8'h00}, /* 0x1318 */
            {8'h00}, /* 0x1317 */
            {8'h00}, /* 0x1316 */
            {8'h00}, /* 0x1315 */
            {8'h00}, /* 0x1314 */
            {8'h00}, /* 0x1313 */
            {8'h00}, /* 0x1312 */
            {8'h00}, /* 0x1311 */
            {8'h00}, /* 0x1310 */
            {8'h00}, /* 0x130f */
            {8'h00}, /* 0x130e */
            {8'h00}, /* 0x130d */
            {8'h00}, /* 0x130c */
            {8'h00}, /* 0x130b */
            {8'h00}, /* 0x130a */
            {8'h00}, /* 0x1309 */
            {8'h00}, /* 0x1308 */
            {8'h00}, /* 0x1307 */
            {8'h00}, /* 0x1306 */
            {8'h00}, /* 0x1305 */
            {8'h00}, /* 0x1304 */
            {8'h00}, /* 0x1303 */
            {8'h00}, /* 0x1302 */
            {8'h00}, /* 0x1301 */
            {8'h00}, /* 0x1300 */
            {8'h00}, /* 0x12ff */
            {8'h00}, /* 0x12fe */
            {8'h00}, /* 0x12fd */
            {8'h00}, /* 0x12fc */
            {8'h00}, /* 0x12fb */
            {8'h00}, /* 0x12fa */
            {8'h00}, /* 0x12f9 */
            {8'h00}, /* 0x12f8 */
            {8'h00}, /* 0x12f7 */
            {8'h00}, /* 0x12f6 */
            {8'h00}, /* 0x12f5 */
            {8'h00}, /* 0x12f4 */
            {8'h00}, /* 0x12f3 */
            {8'h00}, /* 0x12f2 */
            {8'h00}, /* 0x12f1 */
            {8'h00}, /* 0x12f0 */
            {8'h00}, /* 0x12ef */
            {8'h00}, /* 0x12ee */
            {8'h00}, /* 0x12ed */
            {8'h00}, /* 0x12ec */
            {8'h00}, /* 0x12eb */
            {8'h00}, /* 0x12ea */
            {8'h00}, /* 0x12e9 */
            {8'h00}, /* 0x12e8 */
            {8'h00}, /* 0x12e7 */
            {8'h00}, /* 0x12e6 */
            {8'h00}, /* 0x12e5 */
            {8'h00}, /* 0x12e4 */
            {8'h00}, /* 0x12e3 */
            {8'h00}, /* 0x12e2 */
            {8'h00}, /* 0x12e1 */
            {8'h00}, /* 0x12e0 */
            {8'h00}, /* 0x12df */
            {8'h00}, /* 0x12de */
            {8'h00}, /* 0x12dd */
            {8'h00}, /* 0x12dc */
            {8'h00}, /* 0x12db */
            {8'h00}, /* 0x12da */
            {8'h00}, /* 0x12d9 */
            {8'h00}, /* 0x12d8 */
            {8'h00}, /* 0x12d7 */
            {8'h00}, /* 0x12d6 */
            {8'h00}, /* 0x12d5 */
            {8'h00}, /* 0x12d4 */
            {8'h00}, /* 0x12d3 */
            {8'h00}, /* 0x12d2 */
            {8'h00}, /* 0x12d1 */
            {8'h00}, /* 0x12d0 */
            {8'h00}, /* 0x12cf */
            {8'h00}, /* 0x12ce */
            {8'h00}, /* 0x12cd */
            {8'h00}, /* 0x12cc */
            {8'h00}, /* 0x12cb */
            {8'h00}, /* 0x12ca */
            {8'h00}, /* 0x12c9 */
            {8'h00}, /* 0x12c8 */
            {8'h00}, /* 0x12c7 */
            {8'h00}, /* 0x12c6 */
            {8'h00}, /* 0x12c5 */
            {8'h00}, /* 0x12c4 */
            {8'h00}, /* 0x12c3 */
            {8'h00}, /* 0x12c2 */
            {8'h00}, /* 0x12c1 */
            {8'h00}, /* 0x12c0 */
            {8'h00}, /* 0x12bf */
            {8'h00}, /* 0x12be */
            {8'h00}, /* 0x12bd */
            {8'h00}, /* 0x12bc */
            {8'h00}, /* 0x12bb */
            {8'h00}, /* 0x12ba */
            {8'h00}, /* 0x12b9 */
            {8'h00}, /* 0x12b8 */
            {8'h00}, /* 0x12b7 */
            {8'h00}, /* 0x12b6 */
            {8'h00}, /* 0x12b5 */
            {8'h00}, /* 0x12b4 */
            {8'h00}, /* 0x12b3 */
            {8'h00}, /* 0x12b2 */
            {8'h00}, /* 0x12b1 */
            {8'h00}, /* 0x12b0 */
            {8'h00}, /* 0x12af */
            {8'h00}, /* 0x12ae */
            {8'h00}, /* 0x12ad */
            {8'h00}, /* 0x12ac */
            {8'h00}, /* 0x12ab */
            {8'h00}, /* 0x12aa */
            {8'h00}, /* 0x12a9 */
            {8'h00}, /* 0x12a8 */
            {8'h00}, /* 0x12a7 */
            {8'h00}, /* 0x12a6 */
            {8'h00}, /* 0x12a5 */
            {8'h00}, /* 0x12a4 */
            {8'h00}, /* 0x12a3 */
            {8'h00}, /* 0x12a2 */
            {8'h00}, /* 0x12a1 */
            {8'h00}, /* 0x12a0 */
            {8'h00}, /* 0x129f */
            {8'h00}, /* 0x129e */
            {8'h00}, /* 0x129d */
            {8'h00}, /* 0x129c */
            {8'h00}, /* 0x129b */
            {8'h00}, /* 0x129a */
            {8'h00}, /* 0x1299 */
            {8'h00}, /* 0x1298 */
            {8'h00}, /* 0x1297 */
            {8'h00}, /* 0x1296 */
            {8'h00}, /* 0x1295 */
            {8'h00}, /* 0x1294 */
            {8'h00}, /* 0x1293 */
            {8'h00}, /* 0x1292 */
            {8'h00}, /* 0x1291 */
            {8'h00}, /* 0x1290 */
            {8'h00}, /* 0x128f */
            {8'h00}, /* 0x128e */
            {8'h00}, /* 0x128d */
            {8'h00}, /* 0x128c */
            {8'h00}, /* 0x128b */
            {8'h00}, /* 0x128a */
            {8'h00}, /* 0x1289 */
            {8'h00}, /* 0x1288 */
            {8'h00}, /* 0x1287 */
            {8'h00}, /* 0x1286 */
            {8'h00}, /* 0x1285 */
            {8'h00}, /* 0x1284 */
            {8'h00}, /* 0x1283 */
            {8'h00}, /* 0x1282 */
            {8'h00}, /* 0x1281 */
            {8'h00}, /* 0x1280 */
            {8'h00}, /* 0x127f */
            {8'h00}, /* 0x127e */
            {8'h00}, /* 0x127d */
            {8'h00}, /* 0x127c */
            {8'h00}, /* 0x127b */
            {8'h00}, /* 0x127a */
            {8'h00}, /* 0x1279 */
            {8'h00}, /* 0x1278 */
            {8'h00}, /* 0x1277 */
            {8'h00}, /* 0x1276 */
            {8'h00}, /* 0x1275 */
            {8'h00}, /* 0x1274 */
            {8'h00}, /* 0x1273 */
            {8'h00}, /* 0x1272 */
            {8'h00}, /* 0x1271 */
            {8'h00}, /* 0x1270 */
            {8'h00}, /* 0x126f */
            {8'h00}, /* 0x126e */
            {8'h00}, /* 0x126d */
            {8'h00}, /* 0x126c */
            {8'h00}, /* 0x126b */
            {8'h00}, /* 0x126a */
            {8'h00}, /* 0x1269 */
            {8'h00}, /* 0x1268 */
            {8'h00}, /* 0x1267 */
            {8'h00}, /* 0x1266 */
            {8'h00}, /* 0x1265 */
            {8'h00}, /* 0x1264 */
            {8'h00}, /* 0x1263 */
            {8'h00}, /* 0x1262 */
            {8'h00}, /* 0x1261 */
            {8'h00}, /* 0x1260 */
            {8'h00}, /* 0x125f */
            {8'h00}, /* 0x125e */
            {8'h00}, /* 0x125d */
            {8'h00}, /* 0x125c */
            {8'h00}, /* 0x125b */
            {8'h00}, /* 0x125a */
            {8'h00}, /* 0x1259 */
            {8'h00}, /* 0x1258 */
            {8'h00}, /* 0x1257 */
            {8'h00}, /* 0x1256 */
            {8'h00}, /* 0x1255 */
            {8'h00}, /* 0x1254 */
            {8'h00}, /* 0x1253 */
            {8'h00}, /* 0x1252 */
            {8'h00}, /* 0x1251 */
            {8'h00}, /* 0x1250 */
            {8'h00}, /* 0x124f */
            {8'h00}, /* 0x124e */
            {8'h00}, /* 0x124d */
            {8'h00}, /* 0x124c */
            {8'h00}, /* 0x124b */
            {8'h00}, /* 0x124a */
            {8'h00}, /* 0x1249 */
            {8'h00}, /* 0x1248 */
            {8'h00}, /* 0x1247 */
            {8'h00}, /* 0x1246 */
            {8'h00}, /* 0x1245 */
            {8'h00}, /* 0x1244 */
            {8'h00}, /* 0x1243 */
            {8'h00}, /* 0x1242 */
            {8'h00}, /* 0x1241 */
            {8'h00}, /* 0x1240 */
            {8'h00}, /* 0x123f */
            {8'h00}, /* 0x123e */
            {8'h00}, /* 0x123d */
            {8'h00}, /* 0x123c */
            {8'h00}, /* 0x123b */
            {8'h00}, /* 0x123a */
            {8'h00}, /* 0x1239 */
            {8'h00}, /* 0x1238 */
            {8'h00}, /* 0x1237 */
            {8'h00}, /* 0x1236 */
            {8'h00}, /* 0x1235 */
            {8'h00}, /* 0x1234 */
            {8'h00}, /* 0x1233 */
            {8'h00}, /* 0x1232 */
            {8'h00}, /* 0x1231 */
            {8'h00}, /* 0x1230 */
            {8'h00}, /* 0x122f */
            {8'h00}, /* 0x122e */
            {8'h00}, /* 0x122d */
            {8'h00}, /* 0x122c */
            {8'h00}, /* 0x122b */
            {8'h00}, /* 0x122a */
            {8'h00}, /* 0x1229 */
            {8'h00}, /* 0x1228 */
            {8'h00}, /* 0x1227 */
            {8'h00}, /* 0x1226 */
            {8'h00}, /* 0x1225 */
            {8'h00}, /* 0x1224 */
            {8'h00}, /* 0x1223 */
            {8'h00}, /* 0x1222 */
            {8'h00}, /* 0x1221 */
            {8'h00}, /* 0x1220 */
            {8'h00}, /* 0x121f */
            {8'h00}, /* 0x121e */
            {8'h00}, /* 0x121d */
            {8'h00}, /* 0x121c */
            {8'h00}, /* 0x121b */
            {8'h00}, /* 0x121a */
            {8'h00}, /* 0x1219 */
            {8'h00}, /* 0x1218 */
            {8'h00}, /* 0x1217 */
            {8'h00}, /* 0x1216 */
            {8'h00}, /* 0x1215 */
            {8'h00}, /* 0x1214 */
            {8'h00}, /* 0x1213 */
            {8'h00}, /* 0x1212 */
            {8'h00}, /* 0x1211 */
            {8'h00}, /* 0x1210 */
            {8'h00}, /* 0x120f */
            {8'h00}, /* 0x120e */
            {8'h00}, /* 0x120d */
            {8'h00}, /* 0x120c */
            {8'h00}, /* 0x120b */
            {8'h00}, /* 0x120a */
            {8'h00}, /* 0x1209 */
            {8'h00}, /* 0x1208 */
            {8'h00}, /* 0x1207 */
            {8'h00}, /* 0x1206 */
            {8'h00}, /* 0x1205 */
            {8'h00}, /* 0x1204 */
            {8'h00}, /* 0x1203 */
            {8'h00}, /* 0x1202 */
            {8'h00}, /* 0x1201 */
            {8'h00}, /* 0x1200 */
            {8'h00}, /* 0x11ff */
            {8'h00}, /* 0x11fe */
            {8'h00}, /* 0x11fd */
            {8'h00}, /* 0x11fc */
            {8'h00}, /* 0x11fb */
            {8'h00}, /* 0x11fa */
            {8'h00}, /* 0x11f9 */
            {8'h00}, /* 0x11f8 */
            {8'h00}, /* 0x11f7 */
            {8'h00}, /* 0x11f6 */
            {8'h00}, /* 0x11f5 */
            {8'h00}, /* 0x11f4 */
            {8'h00}, /* 0x11f3 */
            {8'h00}, /* 0x11f2 */
            {8'h00}, /* 0x11f1 */
            {8'h00}, /* 0x11f0 */
            {8'h00}, /* 0x11ef */
            {8'h00}, /* 0x11ee */
            {8'h00}, /* 0x11ed */
            {8'h00}, /* 0x11ec */
            {8'h00}, /* 0x11eb */
            {8'h00}, /* 0x11ea */
            {8'h00}, /* 0x11e9 */
            {8'h00}, /* 0x11e8 */
            {8'h00}, /* 0x11e7 */
            {8'h00}, /* 0x11e6 */
            {8'h00}, /* 0x11e5 */
            {8'h00}, /* 0x11e4 */
            {8'h00}, /* 0x11e3 */
            {8'h00}, /* 0x11e2 */
            {8'h00}, /* 0x11e1 */
            {8'h00}, /* 0x11e0 */
            {8'h00}, /* 0x11df */
            {8'h00}, /* 0x11de */
            {8'h00}, /* 0x11dd */
            {8'h00}, /* 0x11dc */
            {8'h00}, /* 0x11db */
            {8'h00}, /* 0x11da */
            {8'h00}, /* 0x11d9 */
            {8'h00}, /* 0x11d8 */
            {8'h00}, /* 0x11d7 */
            {8'h00}, /* 0x11d6 */
            {8'h00}, /* 0x11d5 */
            {8'h00}, /* 0x11d4 */
            {8'h00}, /* 0x11d3 */
            {8'h00}, /* 0x11d2 */
            {8'h00}, /* 0x11d1 */
            {8'h00}, /* 0x11d0 */
            {8'h00}, /* 0x11cf */
            {8'h00}, /* 0x11ce */
            {8'h00}, /* 0x11cd */
            {8'h00}, /* 0x11cc */
            {8'h00}, /* 0x11cb */
            {8'h00}, /* 0x11ca */
            {8'h00}, /* 0x11c9 */
            {8'h00}, /* 0x11c8 */
            {8'h00}, /* 0x11c7 */
            {8'h00}, /* 0x11c6 */
            {8'h00}, /* 0x11c5 */
            {8'h00}, /* 0x11c4 */
            {8'h00}, /* 0x11c3 */
            {8'h00}, /* 0x11c2 */
            {8'h00}, /* 0x11c1 */
            {8'h00}, /* 0x11c0 */
            {8'h00}, /* 0x11bf */
            {8'h00}, /* 0x11be */
            {8'h00}, /* 0x11bd */
            {8'h00}, /* 0x11bc */
            {8'h00}, /* 0x11bb */
            {8'h00}, /* 0x11ba */
            {8'h00}, /* 0x11b9 */
            {8'h00}, /* 0x11b8 */
            {8'h00}, /* 0x11b7 */
            {8'h00}, /* 0x11b6 */
            {8'h00}, /* 0x11b5 */
            {8'h00}, /* 0x11b4 */
            {8'h00}, /* 0x11b3 */
            {8'h00}, /* 0x11b2 */
            {8'h00}, /* 0x11b1 */
            {8'h00}, /* 0x11b0 */
            {8'h00}, /* 0x11af */
            {8'h00}, /* 0x11ae */
            {8'h00}, /* 0x11ad */
            {8'h00}, /* 0x11ac */
            {8'h00}, /* 0x11ab */
            {8'h00}, /* 0x11aa */
            {8'h00}, /* 0x11a9 */
            {8'h00}, /* 0x11a8 */
            {8'h00}, /* 0x11a7 */
            {8'h00}, /* 0x11a6 */
            {8'h00}, /* 0x11a5 */
            {8'h00}, /* 0x11a4 */
            {8'h00}, /* 0x11a3 */
            {8'h00}, /* 0x11a2 */
            {8'h00}, /* 0x11a1 */
            {8'h00}, /* 0x11a0 */
            {8'h00}, /* 0x119f */
            {8'h00}, /* 0x119e */
            {8'h00}, /* 0x119d */
            {8'h00}, /* 0x119c */
            {8'h00}, /* 0x119b */
            {8'h00}, /* 0x119a */
            {8'h00}, /* 0x1199 */
            {8'h00}, /* 0x1198 */
            {8'h00}, /* 0x1197 */
            {8'h00}, /* 0x1196 */
            {8'h00}, /* 0x1195 */
            {8'h00}, /* 0x1194 */
            {8'h00}, /* 0x1193 */
            {8'h00}, /* 0x1192 */
            {8'h00}, /* 0x1191 */
            {8'h00}, /* 0x1190 */
            {8'h00}, /* 0x118f */
            {8'h00}, /* 0x118e */
            {8'h00}, /* 0x118d */
            {8'h00}, /* 0x118c */
            {8'h00}, /* 0x118b */
            {8'h00}, /* 0x118a */
            {8'h00}, /* 0x1189 */
            {8'h00}, /* 0x1188 */
            {8'h00}, /* 0x1187 */
            {8'h00}, /* 0x1186 */
            {8'h00}, /* 0x1185 */
            {8'h00}, /* 0x1184 */
            {8'h00}, /* 0x1183 */
            {8'h00}, /* 0x1182 */
            {8'h00}, /* 0x1181 */
            {8'h00}, /* 0x1180 */
            {8'h00}, /* 0x117f */
            {8'h00}, /* 0x117e */
            {8'h00}, /* 0x117d */
            {8'h00}, /* 0x117c */
            {8'h00}, /* 0x117b */
            {8'h00}, /* 0x117a */
            {8'h00}, /* 0x1179 */
            {8'h00}, /* 0x1178 */
            {8'h00}, /* 0x1177 */
            {8'h00}, /* 0x1176 */
            {8'h00}, /* 0x1175 */
            {8'h00}, /* 0x1174 */
            {8'h00}, /* 0x1173 */
            {8'h00}, /* 0x1172 */
            {8'h00}, /* 0x1171 */
            {8'h00}, /* 0x1170 */
            {8'h00}, /* 0x116f */
            {8'h00}, /* 0x116e */
            {8'h00}, /* 0x116d */
            {8'h00}, /* 0x116c */
            {8'h00}, /* 0x116b */
            {8'h00}, /* 0x116a */
            {8'h00}, /* 0x1169 */
            {8'h00}, /* 0x1168 */
            {8'h00}, /* 0x1167 */
            {8'h00}, /* 0x1166 */
            {8'h00}, /* 0x1165 */
            {8'h00}, /* 0x1164 */
            {8'h00}, /* 0x1163 */
            {8'h00}, /* 0x1162 */
            {8'h00}, /* 0x1161 */
            {8'h00}, /* 0x1160 */
            {8'h00}, /* 0x115f */
            {8'h00}, /* 0x115e */
            {8'h00}, /* 0x115d */
            {8'h00}, /* 0x115c */
            {8'h00}, /* 0x115b */
            {8'h00}, /* 0x115a */
            {8'h00}, /* 0x1159 */
            {8'h00}, /* 0x1158 */
            {8'h00}, /* 0x1157 */
            {8'h00}, /* 0x1156 */
            {8'h00}, /* 0x1155 */
            {8'h00}, /* 0x1154 */
            {8'h00}, /* 0x1153 */
            {8'h00}, /* 0x1152 */
            {8'h00}, /* 0x1151 */
            {8'h00}, /* 0x1150 */
            {8'h00}, /* 0x114f */
            {8'h00}, /* 0x114e */
            {8'h00}, /* 0x114d */
            {8'h00}, /* 0x114c */
            {8'h00}, /* 0x114b */
            {8'h00}, /* 0x114a */
            {8'h00}, /* 0x1149 */
            {8'h00}, /* 0x1148 */
            {8'h00}, /* 0x1147 */
            {8'h00}, /* 0x1146 */
            {8'h00}, /* 0x1145 */
            {8'h00}, /* 0x1144 */
            {8'h00}, /* 0x1143 */
            {8'h00}, /* 0x1142 */
            {8'h00}, /* 0x1141 */
            {8'h00}, /* 0x1140 */
            {8'h00}, /* 0x113f */
            {8'h00}, /* 0x113e */
            {8'h00}, /* 0x113d */
            {8'h00}, /* 0x113c */
            {8'h00}, /* 0x113b */
            {8'h00}, /* 0x113a */
            {8'h00}, /* 0x1139 */
            {8'h00}, /* 0x1138 */
            {8'h00}, /* 0x1137 */
            {8'h00}, /* 0x1136 */
            {8'h00}, /* 0x1135 */
            {8'h00}, /* 0x1134 */
            {8'h00}, /* 0x1133 */
            {8'h00}, /* 0x1132 */
            {8'h00}, /* 0x1131 */
            {8'h00}, /* 0x1130 */
            {8'h00}, /* 0x112f */
            {8'h00}, /* 0x112e */
            {8'h00}, /* 0x112d */
            {8'h00}, /* 0x112c */
            {8'h00}, /* 0x112b */
            {8'h00}, /* 0x112a */
            {8'h00}, /* 0x1129 */
            {8'h00}, /* 0x1128 */
            {8'h00}, /* 0x1127 */
            {8'h00}, /* 0x1126 */
            {8'h00}, /* 0x1125 */
            {8'h00}, /* 0x1124 */
            {8'h00}, /* 0x1123 */
            {8'h00}, /* 0x1122 */
            {8'h00}, /* 0x1121 */
            {8'h00}, /* 0x1120 */
            {8'h00}, /* 0x111f */
            {8'h00}, /* 0x111e */
            {8'h00}, /* 0x111d */
            {8'h00}, /* 0x111c */
            {8'h00}, /* 0x111b */
            {8'h00}, /* 0x111a */
            {8'h00}, /* 0x1119 */
            {8'h00}, /* 0x1118 */
            {8'h00}, /* 0x1117 */
            {8'h00}, /* 0x1116 */
            {8'h00}, /* 0x1115 */
            {8'h00}, /* 0x1114 */
            {8'h00}, /* 0x1113 */
            {8'h00}, /* 0x1112 */
            {8'h00}, /* 0x1111 */
            {8'h00}, /* 0x1110 */
            {8'h00}, /* 0x110f */
            {8'h00}, /* 0x110e */
            {8'h00}, /* 0x110d */
            {8'h00}, /* 0x110c */
            {8'h00}, /* 0x110b */
            {8'h00}, /* 0x110a */
            {8'h00}, /* 0x1109 */
            {8'h00}, /* 0x1108 */
            {8'h00}, /* 0x1107 */
            {8'h00}, /* 0x1106 */
            {8'h00}, /* 0x1105 */
            {8'h00}, /* 0x1104 */
            {8'h00}, /* 0x1103 */
            {8'h00}, /* 0x1102 */
            {8'h00}, /* 0x1101 */
            {8'h00}, /* 0x1100 */
            {8'h00}, /* 0x10ff */
            {8'h00}, /* 0x10fe */
            {8'h00}, /* 0x10fd */
            {8'h00}, /* 0x10fc */
            {8'h00}, /* 0x10fb */
            {8'h00}, /* 0x10fa */
            {8'h00}, /* 0x10f9 */
            {8'h00}, /* 0x10f8 */
            {8'h00}, /* 0x10f7 */
            {8'h00}, /* 0x10f6 */
            {8'h00}, /* 0x10f5 */
            {8'h00}, /* 0x10f4 */
            {8'h00}, /* 0x10f3 */
            {8'h00}, /* 0x10f2 */
            {8'h00}, /* 0x10f1 */
            {8'h00}, /* 0x10f0 */
            {8'h00}, /* 0x10ef */
            {8'h00}, /* 0x10ee */
            {8'h00}, /* 0x10ed */
            {8'h00}, /* 0x10ec */
            {8'h00}, /* 0x10eb */
            {8'h00}, /* 0x10ea */
            {8'h00}, /* 0x10e9 */
            {8'h00}, /* 0x10e8 */
            {8'h00}, /* 0x10e7 */
            {8'h00}, /* 0x10e6 */
            {8'h00}, /* 0x10e5 */
            {8'h00}, /* 0x10e4 */
            {8'h00}, /* 0x10e3 */
            {8'h00}, /* 0x10e2 */
            {8'h00}, /* 0x10e1 */
            {8'h00}, /* 0x10e0 */
            {8'h00}, /* 0x10df */
            {8'h00}, /* 0x10de */
            {8'h00}, /* 0x10dd */
            {8'h00}, /* 0x10dc */
            {8'h00}, /* 0x10db */
            {8'h00}, /* 0x10da */
            {8'h00}, /* 0x10d9 */
            {8'h00}, /* 0x10d8 */
            {8'h00}, /* 0x10d7 */
            {8'h00}, /* 0x10d6 */
            {8'h00}, /* 0x10d5 */
            {8'h00}, /* 0x10d4 */
            {8'h00}, /* 0x10d3 */
            {8'h00}, /* 0x10d2 */
            {8'h00}, /* 0x10d1 */
            {8'h00}, /* 0x10d0 */
            {8'h00}, /* 0x10cf */
            {8'h00}, /* 0x10ce */
            {8'h00}, /* 0x10cd */
            {8'h00}, /* 0x10cc */
            {8'h00}, /* 0x10cb */
            {8'h00}, /* 0x10ca */
            {8'h00}, /* 0x10c9 */
            {8'h00}, /* 0x10c8 */
            {8'h00}, /* 0x10c7 */
            {8'h00}, /* 0x10c6 */
            {8'h00}, /* 0x10c5 */
            {8'h00}, /* 0x10c4 */
            {8'h00}, /* 0x10c3 */
            {8'h00}, /* 0x10c2 */
            {8'h00}, /* 0x10c1 */
            {8'h00}, /* 0x10c0 */
            {8'h00}, /* 0x10bf */
            {8'h00}, /* 0x10be */
            {8'h00}, /* 0x10bd */
            {8'h00}, /* 0x10bc */
            {8'h00}, /* 0x10bb */
            {8'h00}, /* 0x10ba */
            {8'h00}, /* 0x10b9 */
            {8'h00}, /* 0x10b8 */
            {8'h00}, /* 0x10b7 */
            {8'h00}, /* 0x10b6 */
            {8'h00}, /* 0x10b5 */
            {8'h00}, /* 0x10b4 */
            {8'h00}, /* 0x10b3 */
            {8'h00}, /* 0x10b2 */
            {8'h00}, /* 0x10b1 */
            {8'h00}, /* 0x10b0 */
            {8'h00}, /* 0x10af */
            {8'h00}, /* 0x10ae */
            {8'h00}, /* 0x10ad */
            {8'h00}, /* 0x10ac */
            {8'h00}, /* 0x10ab */
            {8'h00}, /* 0x10aa */
            {8'h00}, /* 0x10a9 */
            {8'h00}, /* 0x10a8 */
            {8'h00}, /* 0x10a7 */
            {8'h00}, /* 0x10a6 */
            {8'h00}, /* 0x10a5 */
            {8'h00}, /* 0x10a4 */
            {8'h00}, /* 0x10a3 */
            {8'h00}, /* 0x10a2 */
            {8'h00}, /* 0x10a1 */
            {8'h00}, /* 0x10a0 */
            {8'h00}, /* 0x109f */
            {8'h00}, /* 0x109e */
            {8'h00}, /* 0x109d */
            {8'h00}, /* 0x109c */
            {8'h00}, /* 0x109b */
            {8'h00}, /* 0x109a */
            {8'h00}, /* 0x1099 */
            {8'h00}, /* 0x1098 */
            {8'h00}, /* 0x1097 */
            {8'h00}, /* 0x1096 */
            {8'h00}, /* 0x1095 */
            {8'h00}, /* 0x1094 */
            {8'h00}, /* 0x1093 */
            {8'h00}, /* 0x1092 */
            {8'h00}, /* 0x1091 */
            {8'h00}, /* 0x1090 */
            {8'h00}, /* 0x108f */
            {8'h00}, /* 0x108e */
            {8'h00}, /* 0x108d */
            {8'h00}, /* 0x108c */
            {8'h00}, /* 0x108b */
            {8'h00}, /* 0x108a */
            {8'h00}, /* 0x1089 */
            {8'h00}, /* 0x1088 */
            {8'h00}, /* 0x1087 */
            {8'h00}, /* 0x1086 */
            {8'h00}, /* 0x1085 */
            {8'h00}, /* 0x1084 */
            {8'h00}, /* 0x1083 */
            {8'h00}, /* 0x1082 */
            {8'h00}, /* 0x1081 */
            {8'h00}, /* 0x1080 */
            {8'h00}, /* 0x107f */
            {8'h00}, /* 0x107e */
            {8'h00}, /* 0x107d */
            {8'h00}, /* 0x107c */
            {8'h00}, /* 0x107b */
            {8'h00}, /* 0x107a */
            {8'h00}, /* 0x1079 */
            {8'h00}, /* 0x1078 */
            {8'h00}, /* 0x1077 */
            {8'h00}, /* 0x1076 */
            {8'h00}, /* 0x1075 */
            {8'h00}, /* 0x1074 */
            {8'h00}, /* 0x1073 */
            {8'h00}, /* 0x1072 */
            {8'h00}, /* 0x1071 */
            {8'h00}, /* 0x1070 */
            {8'h00}, /* 0x106f */
            {8'h00}, /* 0x106e */
            {8'h00}, /* 0x106d */
            {8'h00}, /* 0x106c */
            {8'h00}, /* 0x106b */
            {8'h00}, /* 0x106a */
            {8'h00}, /* 0x1069 */
            {8'h00}, /* 0x1068 */
            {8'h00}, /* 0x1067 */
            {8'h00}, /* 0x1066 */
            {8'h00}, /* 0x1065 */
            {8'h00}, /* 0x1064 */
            {8'h00}, /* 0x1063 */
            {8'h00}, /* 0x1062 */
            {8'h00}, /* 0x1061 */
            {8'h00}, /* 0x1060 */
            {8'h00}, /* 0x105f */
            {8'h00}, /* 0x105e */
            {8'h00}, /* 0x105d */
            {8'h00}, /* 0x105c */
            {8'h00}, /* 0x105b */
            {8'h00}, /* 0x105a */
            {8'h00}, /* 0x1059 */
            {8'h00}, /* 0x1058 */
            {8'h00}, /* 0x1057 */
            {8'h00}, /* 0x1056 */
            {8'h00}, /* 0x1055 */
            {8'h00}, /* 0x1054 */
            {8'h00}, /* 0x1053 */
            {8'h00}, /* 0x1052 */
            {8'h00}, /* 0x1051 */
            {8'h00}, /* 0x1050 */
            {8'h00}, /* 0x104f */
            {8'h00}, /* 0x104e */
            {8'h00}, /* 0x104d */
            {8'h00}, /* 0x104c */
            {8'h00}, /* 0x104b */
            {8'h00}, /* 0x104a */
            {8'h00}, /* 0x1049 */
            {8'h00}, /* 0x1048 */
            {8'h00}, /* 0x1047 */
            {8'h00}, /* 0x1046 */
            {8'h00}, /* 0x1045 */
            {8'h00}, /* 0x1044 */
            {8'h00}, /* 0x1043 */
            {8'h00}, /* 0x1042 */
            {8'h00}, /* 0x1041 */
            {8'h00}, /* 0x1040 */
            {8'h00}, /* 0x103f */
            {8'h00}, /* 0x103e */
            {8'h00}, /* 0x103d */
            {8'h00}, /* 0x103c */
            {8'h00}, /* 0x103b */
            {8'h00}, /* 0x103a */
            {8'h00}, /* 0x1039 */
            {8'h00}, /* 0x1038 */
            {8'h00}, /* 0x1037 */
            {8'h00}, /* 0x1036 */
            {8'h00}, /* 0x1035 */
            {8'h00}, /* 0x1034 */
            {8'h00}, /* 0x1033 */
            {8'h00}, /* 0x1032 */
            {8'h00}, /* 0x1031 */
            {8'h00}, /* 0x1030 */
            {8'h00}, /* 0x102f */
            {8'h00}, /* 0x102e */
            {8'h00}, /* 0x102d */
            {8'h00}, /* 0x102c */
            {8'h00}, /* 0x102b */
            {8'h00}, /* 0x102a */
            {8'h00}, /* 0x1029 */
            {8'h00}, /* 0x1028 */
            {8'h00}, /* 0x1027 */
            {8'h00}, /* 0x1026 */
            {8'h00}, /* 0x1025 */
            {8'h00}, /* 0x1024 */
            {8'h00}, /* 0x1023 */
            {8'h00}, /* 0x1022 */
            {8'h00}, /* 0x1021 */
            {8'h00}, /* 0x1020 */
            {8'h00}, /* 0x101f */
            {8'h00}, /* 0x101e */
            {8'h00}, /* 0x101d */
            {8'h00}, /* 0x101c */
            {8'h00}, /* 0x101b */
            {8'h00}, /* 0x101a */
            {8'h00}, /* 0x1019 */
            {8'h00}, /* 0x1018 */
            {8'h00}, /* 0x1017 */
            {8'h00}, /* 0x1016 */
            {8'h00}, /* 0x1015 */
            {8'h00}, /* 0x1014 */
            {8'h00}, /* 0x1013 */
            {8'h00}, /* 0x1012 */
            {8'h00}, /* 0x1011 */
            {8'h00}, /* 0x1010 */
            {8'h00}, /* 0x100f */
            {8'h00}, /* 0x100e */
            {8'h00}, /* 0x100d */
            {8'h00}, /* 0x100c */
            {8'h00}, /* 0x100b */
            {8'h00}, /* 0x100a */
            {8'h00}, /* 0x1009 */
            {8'h00}, /* 0x1008 */
            {8'h00}, /* 0x1007 */
            {8'h00}, /* 0x1006 */
            {8'h00}, /* 0x1005 */
            {8'h00}, /* 0x1004 */
            {8'h00}, /* 0x1003 */
            {8'h00}, /* 0x1002 */
            {8'h00}, /* 0x1001 */
            {8'h00}, /* 0x1000 */
            {8'h00}, /* 0x0fff */
            {8'h00}, /* 0x0ffe */
            {8'h00}, /* 0x0ffd */
            {8'h00}, /* 0x0ffc */
            {8'h00}, /* 0x0ffb */
            {8'h00}, /* 0x0ffa */
            {8'h00}, /* 0x0ff9 */
            {8'h00}, /* 0x0ff8 */
            {8'h00}, /* 0x0ff7 */
            {8'h00}, /* 0x0ff6 */
            {8'h00}, /* 0x0ff5 */
            {8'h00}, /* 0x0ff4 */
            {8'h00}, /* 0x0ff3 */
            {8'h00}, /* 0x0ff2 */
            {8'h00}, /* 0x0ff1 */
            {8'h00}, /* 0x0ff0 */
            {8'h00}, /* 0x0fef */
            {8'h00}, /* 0x0fee */
            {8'h00}, /* 0x0fed */
            {8'h00}, /* 0x0fec */
            {8'h00}, /* 0x0feb */
            {8'h00}, /* 0x0fea */
            {8'h00}, /* 0x0fe9 */
            {8'h00}, /* 0x0fe8 */
            {8'h00}, /* 0x0fe7 */
            {8'h00}, /* 0x0fe6 */
            {8'h00}, /* 0x0fe5 */
            {8'h00}, /* 0x0fe4 */
            {8'h00}, /* 0x0fe3 */
            {8'h00}, /* 0x0fe2 */
            {8'h00}, /* 0x0fe1 */
            {8'h00}, /* 0x0fe0 */
            {8'h00}, /* 0x0fdf */
            {8'h00}, /* 0x0fde */
            {8'h00}, /* 0x0fdd */
            {8'h00}, /* 0x0fdc */
            {8'h00}, /* 0x0fdb */
            {8'h00}, /* 0x0fda */
            {8'h00}, /* 0x0fd9 */
            {8'h00}, /* 0x0fd8 */
            {8'h00}, /* 0x0fd7 */
            {8'h00}, /* 0x0fd6 */
            {8'h00}, /* 0x0fd5 */
            {8'h00}, /* 0x0fd4 */
            {8'h00}, /* 0x0fd3 */
            {8'h00}, /* 0x0fd2 */
            {8'h00}, /* 0x0fd1 */
            {8'h00}, /* 0x0fd0 */
            {8'h00}, /* 0x0fcf */
            {8'h00}, /* 0x0fce */
            {8'h00}, /* 0x0fcd */
            {8'h00}, /* 0x0fcc */
            {8'h00}, /* 0x0fcb */
            {8'h00}, /* 0x0fca */
            {8'h00}, /* 0x0fc9 */
            {8'h00}, /* 0x0fc8 */
            {8'h00}, /* 0x0fc7 */
            {8'h00}, /* 0x0fc6 */
            {8'h00}, /* 0x0fc5 */
            {8'h00}, /* 0x0fc4 */
            {8'h00}, /* 0x0fc3 */
            {8'h00}, /* 0x0fc2 */
            {8'h00}, /* 0x0fc1 */
            {8'h00}, /* 0x0fc0 */
            {8'h00}, /* 0x0fbf */
            {8'h00}, /* 0x0fbe */
            {8'h00}, /* 0x0fbd */
            {8'h00}, /* 0x0fbc */
            {8'h00}, /* 0x0fbb */
            {8'h00}, /* 0x0fba */
            {8'h00}, /* 0x0fb9 */
            {8'h00}, /* 0x0fb8 */
            {8'h00}, /* 0x0fb7 */
            {8'h00}, /* 0x0fb6 */
            {8'h00}, /* 0x0fb5 */
            {8'h00}, /* 0x0fb4 */
            {8'h00}, /* 0x0fb3 */
            {8'h00}, /* 0x0fb2 */
            {8'h00}, /* 0x0fb1 */
            {8'h00}, /* 0x0fb0 */
            {8'h00}, /* 0x0faf */
            {8'h00}, /* 0x0fae */
            {8'h00}, /* 0x0fad */
            {8'h00}, /* 0x0fac */
            {8'h00}, /* 0x0fab */
            {8'h00}, /* 0x0faa */
            {8'h00}, /* 0x0fa9 */
            {8'h00}, /* 0x0fa8 */
            {8'h00}, /* 0x0fa7 */
            {8'h00}, /* 0x0fa6 */
            {8'h00}, /* 0x0fa5 */
            {8'h00}, /* 0x0fa4 */
            {8'h00}, /* 0x0fa3 */
            {8'h00}, /* 0x0fa2 */
            {8'h00}, /* 0x0fa1 */
            {8'h00}, /* 0x0fa0 */
            {8'h00}, /* 0x0f9f */
            {8'h00}, /* 0x0f9e */
            {8'h00}, /* 0x0f9d */
            {8'h00}, /* 0x0f9c */
            {8'h00}, /* 0x0f9b */
            {8'h00}, /* 0x0f9a */
            {8'h00}, /* 0x0f99 */
            {8'h00}, /* 0x0f98 */
            {8'h00}, /* 0x0f97 */
            {8'h00}, /* 0x0f96 */
            {8'h00}, /* 0x0f95 */
            {8'h00}, /* 0x0f94 */
            {8'h00}, /* 0x0f93 */
            {8'h00}, /* 0x0f92 */
            {8'h00}, /* 0x0f91 */
            {8'h00}, /* 0x0f90 */
            {8'h00}, /* 0x0f8f */
            {8'h00}, /* 0x0f8e */
            {8'h00}, /* 0x0f8d */
            {8'h00}, /* 0x0f8c */
            {8'h00}, /* 0x0f8b */
            {8'h00}, /* 0x0f8a */
            {8'h00}, /* 0x0f89 */
            {8'h00}, /* 0x0f88 */
            {8'h00}, /* 0x0f87 */
            {8'h00}, /* 0x0f86 */
            {8'h00}, /* 0x0f85 */
            {8'h00}, /* 0x0f84 */
            {8'h00}, /* 0x0f83 */
            {8'h00}, /* 0x0f82 */
            {8'h00}, /* 0x0f81 */
            {8'h00}, /* 0x0f80 */
            {8'h00}, /* 0x0f7f */
            {8'h00}, /* 0x0f7e */
            {8'h00}, /* 0x0f7d */
            {8'h00}, /* 0x0f7c */
            {8'h00}, /* 0x0f7b */
            {8'h00}, /* 0x0f7a */
            {8'h00}, /* 0x0f79 */
            {8'h00}, /* 0x0f78 */
            {8'h00}, /* 0x0f77 */
            {8'h00}, /* 0x0f76 */
            {8'h00}, /* 0x0f75 */
            {8'h00}, /* 0x0f74 */
            {8'h00}, /* 0x0f73 */
            {8'h00}, /* 0x0f72 */
            {8'h00}, /* 0x0f71 */
            {8'h00}, /* 0x0f70 */
            {8'h00}, /* 0x0f6f */
            {8'h00}, /* 0x0f6e */
            {8'h00}, /* 0x0f6d */
            {8'h00}, /* 0x0f6c */
            {8'h00}, /* 0x0f6b */
            {8'h00}, /* 0x0f6a */
            {8'h00}, /* 0x0f69 */
            {8'h00}, /* 0x0f68 */
            {8'h00}, /* 0x0f67 */
            {8'h00}, /* 0x0f66 */
            {8'h00}, /* 0x0f65 */
            {8'h00}, /* 0x0f64 */
            {8'h00}, /* 0x0f63 */
            {8'h00}, /* 0x0f62 */
            {8'h00}, /* 0x0f61 */
            {8'h00}, /* 0x0f60 */
            {8'h00}, /* 0x0f5f */
            {8'h00}, /* 0x0f5e */
            {8'h00}, /* 0x0f5d */
            {8'h00}, /* 0x0f5c */
            {8'h00}, /* 0x0f5b */
            {8'h00}, /* 0x0f5a */
            {8'h00}, /* 0x0f59 */
            {8'h00}, /* 0x0f58 */
            {8'h00}, /* 0x0f57 */
            {8'h00}, /* 0x0f56 */
            {8'h00}, /* 0x0f55 */
            {8'h00}, /* 0x0f54 */
            {8'h00}, /* 0x0f53 */
            {8'h00}, /* 0x0f52 */
            {8'h00}, /* 0x0f51 */
            {8'h00}, /* 0x0f50 */
            {8'h00}, /* 0x0f4f */
            {8'h00}, /* 0x0f4e */
            {8'h00}, /* 0x0f4d */
            {8'h00}, /* 0x0f4c */
            {8'h00}, /* 0x0f4b */
            {8'h00}, /* 0x0f4a */
            {8'h00}, /* 0x0f49 */
            {8'h00}, /* 0x0f48 */
            {8'h00}, /* 0x0f47 */
            {8'h00}, /* 0x0f46 */
            {8'h00}, /* 0x0f45 */
            {8'h00}, /* 0x0f44 */
            {8'h00}, /* 0x0f43 */
            {8'h00}, /* 0x0f42 */
            {8'h00}, /* 0x0f41 */
            {8'h00}, /* 0x0f40 */
            {8'h00}, /* 0x0f3f */
            {8'h00}, /* 0x0f3e */
            {8'h00}, /* 0x0f3d */
            {8'h00}, /* 0x0f3c */
            {8'h00}, /* 0x0f3b */
            {8'h00}, /* 0x0f3a */
            {8'h00}, /* 0x0f39 */
            {8'h00}, /* 0x0f38 */
            {8'h00}, /* 0x0f37 */
            {8'h00}, /* 0x0f36 */
            {8'h00}, /* 0x0f35 */
            {8'h00}, /* 0x0f34 */
            {8'h00}, /* 0x0f33 */
            {8'h00}, /* 0x0f32 */
            {8'h00}, /* 0x0f31 */
            {8'h00}, /* 0x0f30 */
            {8'h00}, /* 0x0f2f */
            {8'h00}, /* 0x0f2e */
            {8'h00}, /* 0x0f2d */
            {8'h00}, /* 0x0f2c */
            {8'h00}, /* 0x0f2b */
            {8'h00}, /* 0x0f2a */
            {8'h00}, /* 0x0f29 */
            {8'h00}, /* 0x0f28 */
            {8'h00}, /* 0x0f27 */
            {8'h00}, /* 0x0f26 */
            {8'h00}, /* 0x0f25 */
            {8'h00}, /* 0x0f24 */
            {8'h00}, /* 0x0f23 */
            {8'h00}, /* 0x0f22 */
            {8'h00}, /* 0x0f21 */
            {8'h00}, /* 0x0f20 */
            {8'h00}, /* 0x0f1f */
            {8'h00}, /* 0x0f1e */
            {8'h00}, /* 0x0f1d */
            {8'h00}, /* 0x0f1c */
            {8'h00}, /* 0x0f1b */
            {8'h00}, /* 0x0f1a */
            {8'h00}, /* 0x0f19 */
            {8'h00}, /* 0x0f18 */
            {8'h00}, /* 0x0f17 */
            {8'h00}, /* 0x0f16 */
            {8'h00}, /* 0x0f15 */
            {8'h00}, /* 0x0f14 */
            {8'h00}, /* 0x0f13 */
            {8'h00}, /* 0x0f12 */
            {8'h00}, /* 0x0f11 */
            {8'h00}, /* 0x0f10 */
            {8'h00}, /* 0x0f0f */
            {8'h00}, /* 0x0f0e */
            {8'h00}, /* 0x0f0d */
            {8'h00}, /* 0x0f0c */
            {8'h00}, /* 0x0f0b */
            {8'h00}, /* 0x0f0a */
            {8'h00}, /* 0x0f09 */
            {8'h00}, /* 0x0f08 */
            {8'h00}, /* 0x0f07 */
            {8'h00}, /* 0x0f06 */
            {8'h00}, /* 0x0f05 */
            {8'h00}, /* 0x0f04 */
            {8'h00}, /* 0x0f03 */
            {8'h00}, /* 0x0f02 */
            {8'h00}, /* 0x0f01 */
            {8'h00}, /* 0x0f00 */
            {8'h00}, /* 0x0eff */
            {8'h00}, /* 0x0efe */
            {8'h00}, /* 0x0efd */
            {8'h00}, /* 0x0efc */
            {8'h00}, /* 0x0efb */
            {8'h00}, /* 0x0efa */
            {8'h00}, /* 0x0ef9 */
            {8'h00}, /* 0x0ef8 */
            {8'h00}, /* 0x0ef7 */
            {8'h00}, /* 0x0ef6 */
            {8'h00}, /* 0x0ef5 */
            {8'h00}, /* 0x0ef4 */
            {8'h00}, /* 0x0ef3 */
            {8'h00}, /* 0x0ef2 */
            {8'h00}, /* 0x0ef1 */
            {8'h00}, /* 0x0ef0 */
            {8'h00}, /* 0x0eef */
            {8'h00}, /* 0x0eee */
            {8'h00}, /* 0x0eed */
            {8'h00}, /* 0x0eec */
            {8'h00}, /* 0x0eeb */
            {8'h00}, /* 0x0eea */
            {8'h00}, /* 0x0ee9 */
            {8'h00}, /* 0x0ee8 */
            {8'h00}, /* 0x0ee7 */
            {8'h00}, /* 0x0ee6 */
            {8'h00}, /* 0x0ee5 */
            {8'h00}, /* 0x0ee4 */
            {8'h00}, /* 0x0ee3 */
            {8'h00}, /* 0x0ee2 */
            {8'h00}, /* 0x0ee1 */
            {8'h00}, /* 0x0ee0 */
            {8'h00}, /* 0x0edf */
            {8'h00}, /* 0x0ede */
            {8'h00}, /* 0x0edd */
            {8'h00}, /* 0x0edc */
            {8'h00}, /* 0x0edb */
            {8'h00}, /* 0x0eda */
            {8'h00}, /* 0x0ed9 */
            {8'h00}, /* 0x0ed8 */
            {8'h00}, /* 0x0ed7 */
            {8'h00}, /* 0x0ed6 */
            {8'h00}, /* 0x0ed5 */
            {8'h00}, /* 0x0ed4 */
            {8'h00}, /* 0x0ed3 */
            {8'h00}, /* 0x0ed2 */
            {8'h00}, /* 0x0ed1 */
            {8'h00}, /* 0x0ed0 */
            {8'h00}, /* 0x0ecf */
            {8'h00}, /* 0x0ece */
            {8'h00}, /* 0x0ecd */
            {8'h00}, /* 0x0ecc */
            {8'h00}, /* 0x0ecb */
            {8'h00}, /* 0x0eca */
            {8'h00}, /* 0x0ec9 */
            {8'h00}, /* 0x0ec8 */
            {8'h00}, /* 0x0ec7 */
            {8'h00}, /* 0x0ec6 */
            {8'h00}, /* 0x0ec5 */
            {8'h00}, /* 0x0ec4 */
            {8'h00}, /* 0x0ec3 */
            {8'h00}, /* 0x0ec2 */
            {8'h00}, /* 0x0ec1 */
            {8'h00}, /* 0x0ec0 */
            {8'h00}, /* 0x0ebf */
            {8'h00}, /* 0x0ebe */
            {8'h00}, /* 0x0ebd */
            {8'h00}, /* 0x0ebc */
            {8'h00}, /* 0x0ebb */
            {8'h00}, /* 0x0eba */
            {8'h00}, /* 0x0eb9 */
            {8'h00}, /* 0x0eb8 */
            {8'h00}, /* 0x0eb7 */
            {8'h00}, /* 0x0eb6 */
            {8'h00}, /* 0x0eb5 */
            {8'h00}, /* 0x0eb4 */
            {8'h00}, /* 0x0eb3 */
            {8'h00}, /* 0x0eb2 */
            {8'h00}, /* 0x0eb1 */
            {8'h00}, /* 0x0eb0 */
            {8'h00}, /* 0x0eaf */
            {8'h00}, /* 0x0eae */
            {8'h00}, /* 0x0ead */
            {8'h00}, /* 0x0eac */
            {8'h00}, /* 0x0eab */
            {8'h00}, /* 0x0eaa */
            {8'h00}, /* 0x0ea9 */
            {8'h00}, /* 0x0ea8 */
            {8'h00}, /* 0x0ea7 */
            {8'h00}, /* 0x0ea6 */
            {8'h00}, /* 0x0ea5 */
            {8'h00}, /* 0x0ea4 */
            {8'h00}, /* 0x0ea3 */
            {8'h00}, /* 0x0ea2 */
            {8'h00}, /* 0x0ea1 */
            {8'h00}, /* 0x0ea0 */
            {8'h00}, /* 0x0e9f */
            {8'h00}, /* 0x0e9e */
            {8'h00}, /* 0x0e9d */
            {8'h00}, /* 0x0e9c */
            {8'h00}, /* 0x0e9b */
            {8'h00}, /* 0x0e9a */
            {8'h00}, /* 0x0e99 */
            {8'h00}, /* 0x0e98 */
            {8'h00}, /* 0x0e97 */
            {8'h00}, /* 0x0e96 */
            {8'h00}, /* 0x0e95 */
            {8'h00}, /* 0x0e94 */
            {8'h00}, /* 0x0e93 */
            {8'h00}, /* 0x0e92 */
            {8'h00}, /* 0x0e91 */
            {8'h00}, /* 0x0e90 */
            {8'h00}, /* 0x0e8f */
            {8'h00}, /* 0x0e8e */
            {8'h00}, /* 0x0e8d */
            {8'h00}, /* 0x0e8c */
            {8'h00}, /* 0x0e8b */
            {8'h00}, /* 0x0e8a */
            {8'h00}, /* 0x0e89 */
            {8'h00}, /* 0x0e88 */
            {8'h00}, /* 0x0e87 */
            {8'h00}, /* 0x0e86 */
            {8'h00}, /* 0x0e85 */
            {8'h00}, /* 0x0e84 */
            {8'h00}, /* 0x0e83 */
            {8'h00}, /* 0x0e82 */
            {8'h00}, /* 0x0e81 */
            {8'h00}, /* 0x0e80 */
            {8'h00}, /* 0x0e7f */
            {8'h00}, /* 0x0e7e */
            {8'h00}, /* 0x0e7d */
            {8'h00}, /* 0x0e7c */
            {8'h00}, /* 0x0e7b */
            {8'h00}, /* 0x0e7a */
            {8'h00}, /* 0x0e79 */
            {8'h00}, /* 0x0e78 */
            {8'h00}, /* 0x0e77 */
            {8'h00}, /* 0x0e76 */
            {8'h00}, /* 0x0e75 */
            {8'h00}, /* 0x0e74 */
            {8'h00}, /* 0x0e73 */
            {8'h00}, /* 0x0e72 */
            {8'h00}, /* 0x0e71 */
            {8'h00}, /* 0x0e70 */
            {8'h00}, /* 0x0e6f */
            {8'h00}, /* 0x0e6e */
            {8'h00}, /* 0x0e6d */
            {8'h00}, /* 0x0e6c */
            {8'h00}, /* 0x0e6b */
            {8'h00}, /* 0x0e6a */
            {8'h00}, /* 0x0e69 */
            {8'h00}, /* 0x0e68 */
            {8'h00}, /* 0x0e67 */
            {8'h00}, /* 0x0e66 */
            {8'h00}, /* 0x0e65 */
            {8'h00}, /* 0x0e64 */
            {8'h00}, /* 0x0e63 */
            {8'h00}, /* 0x0e62 */
            {8'h00}, /* 0x0e61 */
            {8'h00}, /* 0x0e60 */
            {8'h00}, /* 0x0e5f */
            {8'h00}, /* 0x0e5e */
            {8'h00}, /* 0x0e5d */
            {8'h00}, /* 0x0e5c */
            {8'h00}, /* 0x0e5b */
            {8'h00}, /* 0x0e5a */
            {8'h00}, /* 0x0e59 */
            {8'h00}, /* 0x0e58 */
            {8'h00}, /* 0x0e57 */
            {8'h00}, /* 0x0e56 */
            {8'h00}, /* 0x0e55 */
            {8'h00}, /* 0x0e54 */
            {8'h00}, /* 0x0e53 */
            {8'h00}, /* 0x0e52 */
            {8'h00}, /* 0x0e51 */
            {8'h00}, /* 0x0e50 */
            {8'h00}, /* 0x0e4f */
            {8'h00}, /* 0x0e4e */
            {8'h00}, /* 0x0e4d */
            {8'h00}, /* 0x0e4c */
            {8'h00}, /* 0x0e4b */
            {8'h00}, /* 0x0e4a */
            {8'h00}, /* 0x0e49 */
            {8'h00}, /* 0x0e48 */
            {8'h00}, /* 0x0e47 */
            {8'h00}, /* 0x0e46 */
            {8'h00}, /* 0x0e45 */
            {8'h00}, /* 0x0e44 */
            {8'h00}, /* 0x0e43 */
            {8'h00}, /* 0x0e42 */
            {8'h00}, /* 0x0e41 */
            {8'h00}, /* 0x0e40 */
            {8'h00}, /* 0x0e3f */
            {8'h00}, /* 0x0e3e */
            {8'h00}, /* 0x0e3d */
            {8'h00}, /* 0x0e3c */
            {8'h00}, /* 0x0e3b */
            {8'h00}, /* 0x0e3a */
            {8'h00}, /* 0x0e39 */
            {8'h00}, /* 0x0e38 */
            {8'h00}, /* 0x0e37 */
            {8'h00}, /* 0x0e36 */
            {8'h00}, /* 0x0e35 */
            {8'h00}, /* 0x0e34 */
            {8'h00}, /* 0x0e33 */
            {8'h00}, /* 0x0e32 */
            {8'h00}, /* 0x0e31 */
            {8'h00}, /* 0x0e30 */
            {8'h00}, /* 0x0e2f */
            {8'h00}, /* 0x0e2e */
            {8'h00}, /* 0x0e2d */
            {8'h00}, /* 0x0e2c */
            {8'h00}, /* 0x0e2b */
            {8'h00}, /* 0x0e2a */
            {8'h00}, /* 0x0e29 */
            {8'h00}, /* 0x0e28 */
            {8'h00}, /* 0x0e27 */
            {8'h00}, /* 0x0e26 */
            {8'h00}, /* 0x0e25 */
            {8'h00}, /* 0x0e24 */
            {8'h00}, /* 0x0e23 */
            {8'h00}, /* 0x0e22 */
            {8'h00}, /* 0x0e21 */
            {8'h00}, /* 0x0e20 */
            {8'h00}, /* 0x0e1f */
            {8'h00}, /* 0x0e1e */
            {8'h00}, /* 0x0e1d */
            {8'h00}, /* 0x0e1c */
            {8'h00}, /* 0x0e1b */
            {8'h00}, /* 0x0e1a */
            {8'h00}, /* 0x0e19 */
            {8'h00}, /* 0x0e18 */
            {8'h00}, /* 0x0e17 */
            {8'h00}, /* 0x0e16 */
            {8'h00}, /* 0x0e15 */
            {8'h00}, /* 0x0e14 */
            {8'h00}, /* 0x0e13 */
            {8'h00}, /* 0x0e12 */
            {8'h00}, /* 0x0e11 */
            {8'h00}, /* 0x0e10 */
            {8'h00}, /* 0x0e0f */
            {8'h00}, /* 0x0e0e */
            {8'h00}, /* 0x0e0d */
            {8'h00}, /* 0x0e0c */
            {8'h00}, /* 0x0e0b */
            {8'h00}, /* 0x0e0a */
            {8'h00}, /* 0x0e09 */
            {8'h00}, /* 0x0e08 */
            {8'h00}, /* 0x0e07 */
            {8'h00}, /* 0x0e06 */
            {8'h00}, /* 0x0e05 */
            {8'h00}, /* 0x0e04 */
            {8'h00}, /* 0x0e03 */
            {8'h00}, /* 0x0e02 */
            {8'h00}, /* 0x0e01 */
            {8'h00}, /* 0x0e00 */
            {8'h00}, /* 0x0dff */
            {8'h00}, /* 0x0dfe */
            {8'h00}, /* 0x0dfd */
            {8'h00}, /* 0x0dfc */
            {8'h00}, /* 0x0dfb */
            {8'h00}, /* 0x0dfa */
            {8'h00}, /* 0x0df9 */
            {8'h00}, /* 0x0df8 */
            {8'h00}, /* 0x0df7 */
            {8'h00}, /* 0x0df6 */
            {8'h00}, /* 0x0df5 */
            {8'h00}, /* 0x0df4 */
            {8'h00}, /* 0x0df3 */
            {8'h00}, /* 0x0df2 */
            {8'h00}, /* 0x0df1 */
            {8'h00}, /* 0x0df0 */
            {8'h00}, /* 0x0def */
            {8'h00}, /* 0x0dee */
            {8'h00}, /* 0x0ded */
            {8'h00}, /* 0x0dec */
            {8'h00}, /* 0x0deb */
            {8'h00}, /* 0x0dea */
            {8'h00}, /* 0x0de9 */
            {8'h00}, /* 0x0de8 */
            {8'h00}, /* 0x0de7 */
            {8'h00}, /* 0x0de6 */
            {8'h00}, /* 0x0de5 */
            {8'h00}, /* 0x0de4 */
            {8'h00}, /* 0x0de3 */
            {8'h00}, /* 0x0de2 */
            {8'h00}, /* 0x0de1 */
            {8'h00}, /* 0x0de0 */
            {8'h00}, /* 0x0ddf */
            {8'h00}, /* 0x0dde */
            {8'h00}, /* 0x0ddd */
            {8'h00}, /* 0x0ddc */
            {8'h00}, /* 0x0ddb */
            {8'h00}, /* 0x0dda */
            {8'h00}, /* 0x0dd9 */
            {8'h00}, /* 0x0dd8 */
            {8'h00}, /* 0x0dd7 */
            {8'h00}, /* 0x0dd6 */
            {8'h00}, /* 0x0dd5 */
            {8'h00}, /* 0x0dd4 */
            {8'h00}, /* 0x0dd3 */
            {8'h00}, /* 0x0dd2 */
            {8'h00}, /* 0x0dd1 */
            {8'h00}, /* 0x0dd0 */
            {8'h00}, /* 0x0dcf */
            {8'h00}, /* 0x0dce */
            {8'h00}, /* 0x0dcd */
            {8'h00}, /* 0x0dcc */
            {8'h00}, /* 0x0dcb */
            {8'h00}, /* 0x0dca */
            {8'h00}, /* 0x0dc9 */
            {8'h00}, /* 0x0dc8 */
            {8'h00}, /* 0x0dc7 */
            {8'h00}, /* 0x0dc6 */
            {8'h00}, /* 0x0dc5 */
            {8'h00}, /* 0x0dc4 */
            {8'h00}, /* 0x0dc3 */
            {8'h00}, /* 0x0dc2 */
            {8'h00}, /* 0x0dc1 */
            {8'h00}, /* 0x0dc0 */
            {8'h00}, /* 0x0dbf */
            {8'h00}, /* 0x0dbe */
            {8'h00}, /* 0x0dbd */
            {8'h00}, /* 0x0dbc */
            {8'h00}, /* 0x0dbb */
            {8'h00}, /* 0x0dba */
            {8'h00}, /* 0x0db9 */
            {8'h00}, /* 0x0db8 */
            {8'h00}, /* 0x0db7 */
            {8'h00}, /* 0x0db6 */
            {8'h00}, /* 0x0db5 */
            {8'h00}, /* 0x0db4 */
            {8'h00}, /* 0x0db3 */
            {8'h00}, /* 0x0db2 */
            {8'h00}, /* 0x0db1 */
            {8'h00}, /* 0x0db0 */
            {8'h00}, /* 0x0daf */
            {8'h00}, /* 0x0dae */
            {8'h00}, /* 0x0dad */
            {8'h00}, /* 0x0dac */
            {8'h00}, /* 0x0dab */
            {8'h00}, /* 0x0daa */
            {8'h00}, /* 0x0da9 */
            {8'h00}, /* 0x0da8 */
            {8'h00}, /* 0x0da7 */
            {8'h00}, /* 0x0da6 */
            {8'h00}, /* 0x0da5 */
            {8'h00}, /* 0x0da4 */
            {8'h00}, /* 0x0da3 */
            {8'h00}, /* 0x0da2 */
            {8'h00}, /* 0x0da1 */
            {8'h00}, /* 0x0da0 */
            {8'h00}, /* 0x0d9f */
            {8'h00}, /* 0x0d9e */
            {8'h00}, /* 0x0d9d */
            {8'h00}, /* 0x0d9c */
            {8'h00}, /* 0x0d9b */
            {8'h00}, /* 0x0d9a */
            {8'h00}, /* 0x0d99 */
            {8'h00}, /* 0x0d98 */
            {8'h00}, /* 0x0d97 */
            {8'h00}, /* 0x0d96 */
            {8'h00}, /* 0x0d95 */
            {8'h00}, /* 0x0d94 */
            {8'h00}, /* 0x0d93 */
            {8'h00}, /* 0x0d92 */
            {8'h00}, /* 0x0d91 */
            {8'h00}, /* 0x0d90 */
            {8'h00}, /* 0x0d8f */
            {8'h00}, /* 0x0d8e */
            {8'h00}, /* 0x0d8d */
            {8'h00}, /* 0x0d8c */
            {8'h00}, /* 0x0d8b */
            {8'h00}, /* 0x0d8a */
            {8'h00}, /* 0x0d89 */
            {8'h00}, /* 0x0d88 */
            {8'h00}, /* 0x0d87 */
            {8'h00}, /* 0x0d86 */
            {8'h00}, /* 0x0d85 */
            {8'h00}, /* 0x0d84 */
            {8'h00}, /* 0x0d83 */
            {8'h00}, /* 0x0d82 */
            {8'h00}, /* 0x0d81 */
            {8'h00}, /* 0x0d80 */
            {8'h00}, /* 0x0d7f */
            {8'h00}, /* 0x0d7e */
            {8'h00}, /* 0x0d7d */
            {8'h00}, /* 0x0d7c */
            {8'h00}, /* 0x0d7b */
            {8'h00}, /* 0x0d7a */
            {8'h00}, /* 0x0d79 */
            {8'h00}, /* 0x0d78 */
            {8'h00}, /* 0x0d77 */
            {8'h00}, /* 0x0d76 */
            {8'h00}, /* 0x0d75 */
            {8'h00}, /* 0x0d74 */
            {8'h00}, /* 0x0d73 */
            {8'h00}, /* 0x0d72 */
            {8'h00}, /* 0x0d71 */
            {8'h00}, /* 0x0d70 */
            {8'h00}, /* 0x0d6f */
            {8'h00}, /* 0x0d6e */
            {8'h00}, /* 0x0d6d */
            {8'h00}, /* 0x0d6c */
            {8'h00}, /* 0x0d6b */
            {8'h00}, /* 0x0d6a */
            {8'h00}, /* 0x0d69 */
            {8'h00}, /* 0x0d68 */
            {8'h00}, /* 0x0d67 */
            {8'h00}, /* 0x0d66 */
            {8'h00}, /* 0x0d65 */
            {8'h00}, /* 0x0d64 */
            {8'h00}, /* 0x0d63 */
            {8'h00}, /* 0x0d62 */
            {8'h00}, /* 0x0d61 */
            {8'h00}, /* 0x0d60 */
            {8'h00}, /* 0x0d5f */
            {8'h00}, /* 0x0d5e */
            {8'h00}, /* 0x0d5d */
            {8'h00}, /* 0x0d5c */
            {8'h00}, /* 0x0d5b */
            {8'h00}, /* 0x0d5a */
            {8'h00}, /* 0x0d59 */
            {8'h00}, /* 0x0d58 */
            {8'h00}, /* 0x0d57 */
            {8'h00}, /* 0x0d56 */
            {8'h00}, /* 0x0d55 */
            {8'h00}, /* 0x0d54 */
            {8'h00}, /* 0x0d53 */
            {8'h00}, /* 0x0d52 */
            {8'h00}, /* 0x0d51 */
            {8'h00}, /* 0x0d50 */
            {8'h00}, /* 0x0d4f */
            {8'h00}, /* 0x0d4e */
            {8'h00}, /* 0x0d4d */
            {8'h00}, /* 0x0d4c */
            {8'h00}, /* 0x0d4b */
            {8'h00}, /* 0x0d4a */
            {8'h00}, /* 0x0d49 */
            {8'h00}, /* 0x0d48 */
            {8'h00}, /* 0x0d47 */
            {8'h00}, /* 0x0d46 */
            {8'h00}, /* 0x0d45 */
            {8'h00}, /* 0x0d44 */
            {8'h00}, /* 0x0d43 */
            {8'h00}, /* 0x0d42 */
            {8'h00}, /* 0x0d41 */
            {8'h00}, /* 0x0d40 */
            {8'h00}, /* 0x0d3f */
            {8'h00}, /* 0x0d3e */
            {8'h00}, /* 0x0d3d */
            {8'h00}, /* 0x0d3c */
            {8'h00}, /* 0x0d3b */
            {8'h00}, /* 0x0d3a */
            {8'h00}, /* 0x0d39 */
            {8'h00}, /* 0x0d38 */
            {8'h00}, /* 0x0d37 */
            {8'h00}, /* 0x0d36 */
            {8'h00}, /* 0x0d35 */
            {8'h00}, /* 0x0d34 */
            {8'h00}, /* 0x0d33 */
            {8'h00}, /* 0x0d32 */
            {8'h00}, /* 0x0d31 */
            {8'h00}, /* 0x0d30 */
            {8'h00}, /* 0x0d2f */
            {8'h00}, /* 0x0d2e */
            {8'h00}, /* 0x0d2d */
            {8'h00}, /* 0x0d2c */
            {8'h00}, /* 0x0d2b */
            {8'h00}, /* 0x0d2a */
            {8'h00}, /* 0x0d29 */
            {8'h00}, /* 0x0d28 */
            {8'h00}, /* 0x0d27 */
            {8'h00}, /* 0x0d26 */
            {8'h00}, /* 0x0d25 */
            {8'h00}, /* 0x0d24 */
            {8'h00}, /* 0x0d23 */
            {8'h00}, /* 0x0d22 */
            {8'h00}, /* 0x0d21 */
            {8'h00}, /* 0x0d20 */
            {8'h00}, /* 0x0d1f */
            {8'h00}, /* 0x0d1e */
            {8'h00}, /* 0x0d1d */
            {8'h00}, /* 0x0d1c */
            {8'h00}, /* 0x0d1b */
            {8'h00}, /* 0x0d1a */
            {8'h00}, /* 0x0d19 */
            {8'h00}, /* 0x0d18 */
            {8'h00}, /* 0x0d17 */
            {8'h00}, /* 0x0d16 */
            {8'h00}, /* 0x0d15 */
            {8'h00}, /* 0x0d14 */
            {8'h00}, /* 0x0d13 */
            {8'h00}, /* 0x0d12 */
            {8'h00}, /* 0x0d11 */
            {8'h00}, /* 0x0d10 */
            {8'h00}, /* 0x0d0f */
            {8'h00}, /* 0x0d0e */
            {8'h00}, /* 0x0d0d */
            {8'h00}, /* 0x0d0c */
            {8'h00}, /* 0x0d0b */
            {8'h00}, /* 0x0d0a */
            {8'h00}, /* 0x0d09 */
            {8'h00}, /* 0x0d08 */
            {8'h00}, /* 0x0d07 */
            {8'h00}, /* 0x0d06 */
            {8'h00}, /* 0x0d05 */
            {8'h00}, /* 0x0d04 */
            {8'h00}, /* 0x0d03 */
            {8'h00}, /* 0x0d02 */
            {8'h00}, /* 0x0d01 */
            {8'h00}, /* 0x0d00 */
            {8'h00}, /* 0x0cff */
            {8'h00}, /* 0x0cfe */
            {8'h00}, /* 0x0cfd */
            {8'h00}, /* 0x0cfc */
            {8'h00}, /* 0x0cfb */
            {8'h00}, /* 0x0cfa */
            {8'h00}, /* 0x0cf9 */
            {8'h00}, /* 0x0cf8 */
            {8'h00}, /* 0x0cf7 */
            {8'h00}, /* 0x0cf6 */
            {8'h00}, /* 0x0cf5 */
            {8'h00}, /* 0x0cf4 */
            {8'h00}, /* 0x0cf3 */
            {8'h00}, /* 0x0cf2 */
            {8'h00}, /* 0x0cf1 */
            {8'h00}, /* 0x0cf0 */
            {8'h00}, /* 0x0cef */
            {8'h00}, /* 0x0cee */
            {8'h00}, /* 0x0ced */
            {8'h00}, /* 0x0cec */
            {8'h00}, /* 0x0ceb */
            {8'h00}, /* 0x0cea */
            {8'h00}, /* 0x0ce9 */
            {8'h00}, /* 0x0ce8 */
            {8'h00}, /* 0x0ce7 */
            {8'h00}, /* 0x0ce6 */
            {8'h00}, /* 0x0ce5 */
            {8'h00}, /* 0x0ce4 */
            {8'h00}, /* 0x0ce3 */
            {8'h00}, /* 0x0ce2 */
            {8'h00}, /* 0x0ce1 */
            {8'h00}, /* 0x0ce0 */
            {8'h00}, /* 0x0cdf */
            {8'h00}, /* 0x0cde */
            {8'h00}, /* 0x0cdd */
            {8'h00}, /* 0x0cdc */
            {8'h00}, /* 0x0cdb */
            {8'h00}, /* 0x0cda */
            {8'h00}, /* 0x0cd9 */
            {8'h00}, /* 0x0cd8 */
            {8'h00}, /* 0x0cd7 */
            {8'h00}, /* 0x0cd6 */
            {8'h00}, /* 0x0cd5 */
            {8'h00}, /* 0x0cd4 */
            {8'h00}, /* 0x0cd3 */
            {8'h00}, /* 0x0cd2 */
            {8'h00}, /* 0x0cd1 */
            {8'h00}, /* 0x0cd0 */
            {8'h00}, /* 0x0ccf */
            {8'h00}, /* 0x0cce */
            {8'h00}, /* 0x0ccd */
            {8'h00}, /* 0x0ccc */
            {8'h00}, /* 0x0ccb */
            {8'h00}, /* 0x0cca */
            {8'h00}, /* 0x0cc9 */
            {8'h00}, /* 0x0cc8 */
            {8'h00}, /* 0x0cc7 */
            {8'h00}, /* 0x0cc6 */
            {8'h00}, /* 0x0cc5 */
            {8'h00}, /* 0x0cc4 */
            {8'h00}, /* 0x0cc3 */
            {8'h00}, /* 0x0cc2 */
            {8'h00}, /* 0x0cc1 */
            {8'h00}, /* 0x0cc0 */
            {8'h00}, /* 0x0cbf */
            {8'h00}, /* 0x0cbe */
            {8'h00}, /* 0x0cbd */
            {8'h00}, /* 0x0cbc */
            {8'h00}, /* 0x0cbb */
            {8'h00}, /* 0x0cba */
            {8'h00}, /* 0x0cb9 */
            {8'h00}, /* 0x0cb8 */
            {8'h00}, /* 0x0cb7 */
            {8'h00}, /* 0x0cb6 */
            {8'h00}, /* 0x0cb5 */
            {8'h00}, /* 0x0cb4 */
            {8'h00}, /* 0x0cb3 */
            {8'h00}, /* 0x0cb2 */
            {8'h00}, /* 0x0cb1 */
            {8'h00}, /* 0x0cb0 */
            {8'h00}, /* 0x0caf */
            {8'h00}, /* 0x0cae */
            {8'h00}, /* 0x0cad */
            {8'h00}, /* 0x0cac */
            {8'h00}, /* 0x0cab */
            {8'h00}, /* 0x0caa */
            {8'h00}, /* 0x0ca9 */
            {8'h00}, /* 0x0ca8 */
            {8'h00}, /* 0x0ca7 */
            {8'h00}, /* 0x0ca6 */
            {8'h00}, /* 0x0ca5 */
            {8'h00}, /* 0x0ca4 */
            {8'h00}, /* 0x0ca3 */
            {8'h00}, /* 0x0ca2 */
            {8'h00}, /* 0x0ca1 */
            {8'h00}, /* 0x0ca0 */
            {8'h00}, /* 0x0c9f */
            {8'h00}, /* 0x0c9e */
            {8'h00}, /* 0x0c9d */
            {8'h00}, /* 0x0c9c */
            {8'h00}, /* 0x0c9b */
            {8'h00}, /* 0x0c9a */
            {8'h00}, /* 0x0c99 */
            {8'h00}, /* 0x0c98 */
            {8'h00}, /* 0x0c97 */
            {8'h00}, /* 0x0c96 */
            {8'h00}, /* 0x0c95 */
            {8'h00}, /* 0x0c94 */
            {8'h00}, /* 0x0c93 */
            {8'h00}, /* 0x0c92 */
            {8'h00}, /* 0x0c91 */
            {8'h00}, /* 0x0c90 */
            {8'h00}, /* 0x0c8f */
            {8'h00}, /* 0x0c8e */
            {8'h00}, /* 0x0c8d */
            {8'h00}, /* 0x0c8c */
            {8'h00}, /* 0x0c8b */
            {8'h00}, /* 0x0c8a */
            {8'h00}, /* 0x0c89 */
            {8'h00}, /* 0x0c88 */
            {8'h00}, /* 0x0c87 */
            {8'h00}, /* 0x0c86 */
            {8'h00}, /* 0x0c85 */
            {8'h00}, /* 0x0c84 */
            {8'h00}, /* 0x0c83 */
            {8'h00}, /* 0x0c82 */
            {8'h00}, /* 0x0c81 */
            {8'h00}, /* 0x0c80 */
            {8'h00}, /* 0x0c7f */
            {8'h00}, /* 0x0c7e */
            {8'h00}, /* 0x0c7d */
            {8'h00}, /* 0x0c7c */
            {8'h00}, /* 0x0c7b */
            {8'h00}, /* 0x0c7a */
            {8'h00}, /* 0x0c79 */
            {8'h00}, /* 0x0c78 */
            {8'h00}, /* 0x0c77 */
            {8'h00}, /* 0x0c76 */
            {8'h00}, /* 0x0c75 */
            {8'h00}, /* 0x0c74 */
            {8'h00}, /* 0x0c73 */
            {8'h00}, /* 0x0c72 */
            {8'h00}, /* 0x0c71 */
            {8'h00}, /* 0x0c70 */
            {8'h00}, /* 0x0c6f */
            {8'h00}, /* 0x0c6e */
            {8'h00}, /* 0x0c6d */
            {8'h00}, /* 0x0c6c */
            {8'h00}, /* 0x0c6b */
            {8'h00}, /* 0x0c6a */
            {8'h00}, /* 0x0c69 */
            {8'h00}, /* 0x0c68 */
            {8'h00}, /* 0x0c67 */
            {8'h00}, /* 0x0c66 */
            {8'h00}, /* 0x0c65 */
            {8'h00}, /* 0x0c64 */
            {8'h00}, /* 0x0c63 */
            {8'h00}, /* 0x0c62 */
            {8'h00}, /* 0x0c61 */
            {8'h00}, /* 0x0c60 */
            {8'h00}, /* 0x0c5f */
            {8'h00}, /* 0x0c5e */
            {8'h00}, /* 0x0c5d */
            {8'h00}, /* 0x0c5c */
            {8'h00}, /* 0x0c5b */
            {8'h00}, /* 0x0c5a */
            {8'h00}, /* 0x0c59 */
            {8'h00}, /* 0x0c58 */
            {8'h00}, /* 0x0c57 */
            {8'h00}, /* 0x0c56 */
            {8'h00}, /* 0x0c55 */
            {8'h00}, /* 0x0c54 */
            {8'h00}, /* 0x0c53 */
            {8'h00}, /* 0x0c52 */
            {8'h00}, /* 0x0c51 */
            {8'h00}, /* 0x0c50 */
            {8'h00}, /* 0x0c4f */
            {8'h00}, /* 0x0c4e */
            {8'h00}, /* 0x0c4d */
            {8'h00}, /* 0x0c4c */
            {8'h00}, /* 0x0c4b */
            {8'h00}, /* 0x0c4a */
            {8'h00}, /* 0x0c49 */
            {8'h00}, /* 0x0c48 */
            {8'h00}, /* 0x0c47 */
            {8'h00}, /* 0x0c46 */
            {8'h00}, /* 0x0c45 */
            {8'h00}, /* 0x0c44 */
            {8'h00}, /* 0x0c43 */
            {8'h00}, /* 0x0c42 */
            {8'h00}, /* 0x0c41 */
            {8'h00}, /* 0x0c40 */
            {8'h00}, /* 0x0c3f */
            {8'h00}, /* 0x0c3e */
            {8'h00}, /* 0x0c3d */
            {8'h00}, /* 0x0c3c */
            {8'h00}, /* 0x0c3b */
            {8'h00}, /* 0x0c3a */
            {8'h00}, /* 0x0c39 */
            {8'h00}, /* 0x0c38 */
            {8'h00}, /* 0x0c37 */
            {8'h00}, /* 0x0c36 */
            {8'h00}, /* 0x0c35 */
            {8'h00}, /* 0x0c34 */
            {8'h00}, /* 0x0c33 */
            {8'h00}, /* 0x0c32 */
            {8'h00}, /* 0x0c31 */
            {8'h00}, /* 0x0c30 */
            {8'h00}, /* 0x0c2f */
            {8'h00}, /* 0x0c2e */
            {8'h00}, /* 0x0c2d */
            {8'h00}, /* 0x0c2c */
            {8'h00}, /* 0x0c2b */
            {8'h00}, /* 0x0c2a */
            {8'h00}, /* 0x0c29 */
            {8'h00}, /* 0x0c28 */
            {8'h00}, /* 0x0c27 */
            {8'h00}, /* 0x0c26 */
            {8'h00}, /* 0x0c25 */
            {8'h00}, /* 0x0c24 */
            {8'h00}, /* 0x0c23 */
            {8'h00}, /* 0x0c22 */
            {8'h00}, /* 0x0c21 */
            {8'h00}, /* 0x0c20 */
            {8'h00}, /* 0x0c1f */
            {8'h00}, /* 0x0c1e */
            {8'h00}, /* 0x0c1d */
            {8'h00}, /* 0x0c1c */
            {8'h00}, /* 0x0c1b */
            {8'h00}, /* 0x0c1a */
            {8'h00}, /* 0x0c19 */
            {8'h00}, /* 0x0c18 */
            {8'h00}, /* 0x0c17 */
            {8'h00}, /* 0x0c16 */
            {8'h00}, /* 0x0c15 */
            {8'h00}, /* 0x0c14 */
            {8'h00}, /* 0x0c13 */
            {8'h00}, /* 0x0c12 */
            {8'h00}, /* 0x0c11 */
            {8'h00}, /* 0x0c10 */
            {8'h00}, /* 0x0c0f */
            {8'h00}, /* 0x0c0e */
            {8'h00}, /* 0x0c0d */
            {8'h00}, /* 0x0c0c */
            {8'h00}, /* 0x0c0b */
            {8'h00}, /* 0x0c0a */
            {8'h00}, /* 0x0c09 */
            {8'h00}, /* 0x0c08 */
            {8'h00}, /* 0x0c07 */
            {8'h00}, /* 0x0c06 */
            {8'h00}, /* 0x0c05 */
            {8'h00}, /* 0x0c04 */
            {8'h00}, /* 0x0c03 */
            {8'h00}, /* 0x0c02 */
            {8'h00}, /* 0x0c01 */
            {8'h00}, /* 0x0c00 */
            {8'h00}, /* 0x0bff */
            {8'h00}, /* 0x0bfe */
            {8'h00}, /* 0x0bfd */
            {8'h00}, /* 0x0bfc */
            {8'h00}, /* 0x0bfb */
            {8'h00}, /* 0x0bfa */
            {8'h00}, /* 0x0bf9 */
            {8'h00}, /* 0x0bf8 */
            {8'h00}, /* 0x0bf7 */
            {8'h00}, /* 0x0bf6 */
            {8'h00}, /* 0x0bf5 */
            {8'h00}, /* 0x0bf4 */
            {8'h00}, /* 0x0bf3 */
            {8'h00}, /* 0x0bf2 */
            {8'h00}, /* 0x0bf1 */
            {8'h00}, /* 0x0bf0 */
            {8'h00}, /* 0x0bef */
            {8'h00}, /* 0x0bee */
            {8'h00}, /* 0x0bed */
            {8'h00}, /* 0x0bec */
            {8'h00}, /* 0x0beb */
            {8'h00}, /* 0x0bea */
            {8'h00}, /* 0x0be9 */
            {8'h00}, /* 0x0be8 */
            {8'h00}, /* 0x0be7 */
            {8'h00}, /* 0x0be6 */
            {8'h00}, /* 0x0be5 */
            {8'h00}, /* 0x0be4 */
            {8'h00}, /* 0x0be3 */
            {8'h00}, /* 0x0be2 */
            {8'h00}, /* 0x0be1 */
            {8'h00}, /* 0x0be0 */
            {8'h00}, /* 0x0bdf */
            {8'h00}, /* 0x0bde */
            {8'h00}, /* 0x0bdd */
            {8'h00}, /* 0x0bdc */
            {8'h00}, /* 0x0bdb */
            {8'h00}, /* 0x0bda */
            {8'h00}, /* 0x0bd9 */
            {8'h00}, /* 0x0bd8 */
            {8'h00}, /* 0x0bd7 */
            {8'h00}, /* 0x0bd6 */
            {8'h00}, /* 0x0bd5 */
            {8'h00}, /* 0x0bd4 */
            {8'h00}, /* 0x0bd3 */
            {8'h00}, /* 0x0bd2 */
            {8'h00}, /* 0x0bd1 */
            {8'h00}, /* 0x0bd0 */
            {8'h00}, /* 0x0bcf */
            {8'h00}, /* 0x0bce */
            {8'h00}, /* 0x0bcd */
            {8'h00}, /* 0x0bcc */
            {8'h00}, /* 0x0bcb */
            {8'h00}, /* 0x0bca */
            {8'h00}, /* 0x0bc9 */
            {8'h00}, /* 0x0bc8 */
            {8'h00}, /* 0x0bc7 */
            {8'h00}, /* 0x0bc6 */
            {8'h00}, /* 0x0bc5 */
            {8'h00}, /* 0x0bc4 */
            {8'h00}, /* 0x0bc3 */
            {8'h00}, /* 0x0bc2 */
            {8'h00}, /* 0x0bc1 */
            {8'h00}, /* 0x0bc0 */
            {8'h00}, /* 0x0bbf */
            {8'h00}, /* 0x0bbe */
            {8'h00}, /* 0x0bbd */
            {8'h00}, /* 0x0bbc */
            {8'h00}, /* 0x0bbb */
            {8'h00}, /* 0x0bba */
            {8'h00}, /* 0x0bb9 */
            {8'h00}, /* 0x0bb8 */
            {8'h00}, /* 0x0bb7 */
            {8'h00}, /* 0x0bb6 */
            {8'h00}, /* 0x0bb5 */
            {8'h00}, /* 0x0bb4 */
            {8'h00}, /* 0x0bb3 */
            {8'h00}, /* 0x0bb2 */
            {8'h00}, /* 0x0bb1 */
            {8'h00}, /* 0x0bb0 */
            {8'h00}, /* 0x0baf */
            {8'h00}, /* 0x0bae */
            {8'h00}, /* 0x0bad */
            {8'h00}, /* 0x0bac */
            {8'h00}, /* 0x0bab */
            {8'h00}, /* 0x0baa */
            {8'h00}, /* 0x0ba9 */
            {8'h00}, /* 0x0ba8 */
            {8'h00}, /* 0x0ba7 */
            {8'h00}, /* 0x0ba6 */
            {8'h00}, /* 0x0ba5 */
            {8'h00}, /* 0x0ba4 */
            {8'h00}, /* 0x0ba3 */
            {8'h00}, /* 0x0ba2 */
            {8'h00}, /* 0x0ba1 */
            {8'h00}, /* 0x0ba0 */
            {8'h00}, /* 0x0b9f */
            {8'h00}, /* 0x0b9e */
            {8'h00}, /* 0x0b9d */
            {8'h00}, /* 0x0b9c */
            {8'h00}, /* 0x0b9b */
            {8'h00}, /* 0x0b9a */
            {8'h00}, /* 0x0b99 */
            {8'h00}, /* 0x0b98 */
            {8'h00}, /* 0x0b97 */
            {8'h00}, /* 0x0b96 */
            {8'h00}, /* 0x0b95 */
            {8'h00}, /* 0x0b94 */
            {8'h00}, /* 0x0b93 */
            {8'h00}, /* 0x0b92 */
            {8'h00}, /* 0x0b91 */
            {8'h00}, /* 0x0b90 */
            {8'h00}, /* 0x0b8f */
            {8'h00}, /* 0x0b8e */
            {8'h00}, /* 0x0b8d */
            {8'h00}, /* 0x0b8c */
            {8'h00}, /* 0x0b8b */
            {8'h00}, /* 0x0b8a */
            {8'h00}, /* 0x0b89 */
            {8'h00}, /* 0x0b88 */
            {8'h00}, /* 0x0b87 */
            {8'h00}, /* 0x0b86 */
            {8'h00}, /* 0x0b85 */
            {8'h00}, /* 0x0b84 */
            {8'h00}, /* 0x0b83 */
            {8'h00}, /* 0x0b82 */
            {8'h00}, /* 0x0b81 */
            {8'h00}, /* 0x0b80 */
            {8'h00}, /* 0x0b7f */
            {8'h00}, /* 0x0b7e */
            {8'h00}, /* 0x0b7d */
            {8'h00}, /* 0x0b7c */
            {8'h00}, /* 0x0b7b */
            {8'h00}, /* 0x0b7a */
            {8'h00}, /* 0x0b79 */
            {8'h00}, /* 0x0b78 */
            {8'h00}, /* 0x0b77 */
            {8'h00}, /* 0x0b76 */
            {8'h00}, /* 0x0b75 */
            {8'h00}, /* 0x0b74 */
            {8'h00}, /* 0x0b73 */
            {8'h00}, /* 0x0b72 */
            {8'h00}, /* 0x0b71 */
            {8'h00}, /* 0x0b70 */
            {8'h00}, /* 0x0b6f */
            {8'h00}, /* 0x0b6e */
            {8'h00}, /* 0x0b6d */
            {8'h00}, /* 0x0b6c */
            {8'h00}, /* 0x0b6b */
            {8'h00}, /* 0x0b6a */
            {8'h00}, /* 0x0b69 */
            {8'h00}, /* 0x0b68 */
            {8'h00}, /* 0x0b67 */
            {8'h00}, /* 0x0b66 */
            {8'h00}, /* 0x0b65 */
            {8'h00}, /* 0x0b64 */
            {8'h00}, /* 0x0b63 */
            {8'h00}, /* 0x0b62 */
            {8'h00}, /* 0x0b61 */
            {8'h00}, /* 0x0b60 */
            {8'h00}, /* 0x0b5f */
            {8'h00}, /* 0x0b5e */
            {8'h00}, /* 0x0b5d */
            {8'h00}, /* 0x0b5c */
            {8'h00}, /* 0x0b5b */
            {8'h00}, /* 0x0b5a */
            {8'h00}, /* 0x0b59 */
            {8'h00}, /* 0x0b58 */
            {8'h00}, /* 0x0b57 */
            {8'h00}, /* 0x0b56 */
            {8'h00}, /* 0x0b55 */
            {8'h00}, /* 0x0b54 */
            {8'h00}, /* 0x0b53 */
            {8'h00}, /* 0x0b52 */
            {8'h00}, /* 0x0b51 */
            {8'h00}, /* 0x0b50 */
            {8'h00}, /* 0x0b4f */
            {8'h00}, /* 0x0b4e */
            {8'h00}, /* 0x0b4d */
            {8'h00}, /* 0x0b4c */
            {8'h00}, /* 0x0b4b */
            {8'h00}, /* 0x0b4a */
            {8'h00}, /* 0x0b49 */
            {8'h00}, /* 0x0b48 */
            {8'h00}, /* 0x0b47 */
            {8'h00}, /* 0x0b46 */
            {8'h00}, /* 0x0b45 */
            {8'h00}, /* 0x0b44 */
            {8'h00}, /* 0x0b43 */
            {8'h00}, /* 0x0b42 */
            {8'h00}, /* 0x0b41 */
            {8'h00}, /* 0x0b40 */
            {8'h00}, /* 0x0b3f */
            {8'h00}, /* 0x0b3e */
            {8'h00}, /* 0x0b3d */
            {8'h00}, /* 0x0b3c */
            {8'h00}, /* 0x0b3b */
            {8'h00}, /* 0x0b3a */
            {8'h00}, /* 0x0b39 */
            {8'h00}, /* 0x0b38 */
            {8'h00}, /* 0x0b37 */
            {8'h00}, /* 0x0b36 */
            {8'h00}, /* 0x0b35 */
            {8'h00}, /* 0x0b34 */
            {8'h00}, /* 0x0b33 */
            {8'h00}, /* 0x0b32 */
            {8'h00}, /* 0x0b31 */
            {8'h00}, /* 0x0b30 */
            {8'h00}, /* 0x0b2f */
            {8'h00}, /* 0x0b2e */
            {8'h00}, /* 0x0b2d */
            {8'h00}, /* 0x0b2c */
            {8'h00}, /* 0x0b2b */
            {8'h00}, /* 0x0b2a */
            {8'h00}, /* 0x0b29 */
            {8'h00}, /* 0x0b28 */
            {8'h00}, /* 0x0b27 */
            {8'h00}, /* 0x0b26 */
            {8'h00}, /* 0x0b25 */
            {8'h00}, /* 0x0b24 */
            {8'h00}, /* 0x0b23 */
            {8'h00}, /* 0x0b22 */
            {8'h00}, /* 0x0b21 */
            {8'h00}, /* 0x0b20 */
            {8'h00}, /* 0x0b1f */
            {8'h00}, /* 0x0b1e */
            {8'h00}, /* 0x0b1d */
            {8'h00}, /* 0x0b1c */
            {8'h00}, /* 0x0b1b */
            {8'h00}, /* 0x0b1a */
            {8'h00}, /* 0x0b19 */
            {8'h00}, /* 0x0b18 */
            {8'h00}, /* 0x0b17 */
            {8'h00}, /* 0x0b16 */
            {8'h00}, /* 0x0b15 */
            {8'h00}, /* 0x0b14 */
            {8'h00}, /* 0x0b13 */
            {8'h00}, /* 0x0b12 */
            {8'h00}, /* 0x0b11 */
            {8'h00}, /* 0x0b10 */
            {8'h00}, /* 0x0b0f */
            {8'h00}, /* 0x0b0e */
            {8'h00}, /* 0x0b0d */
            {8'h00}, /* 0x0b0c */
            {8'h00}, /* 0x0b0b */
            {8'h00}, /* 0x0b0a */
            {8'h00}, /* 0x0b09 */
            {8'h00}, /* 0x0b08 */
            {8'h00}, /* 0x0b07 */
            {8'h00}, /* 0x0b06 */
            {8'h00}, /* 0x0b05 */
            {8'h00}, /* 0x0b04 */
            {8'h00}, /* 0x0b03 */
            {8'h00}, /* 0x0b02 */
            {8'h00}, /* 0x0b01 */
            {8'h00}, /* 0x0b00 */
            {8'h00}, /* 0x0aff */
            {8'h00}, /* 0x0afe */
            {8'h00}, /* 0x0afd */
            {8'h00}, /* 0x0afc */
            {8'h00}, /* 0x0afb */
            {8'h00}, /* 0x0afa */
            {8'h00}, /* 0x0af9 */
            {8'h00}, /* 0x0af8 */
            {8'h00}, /* 0x0af7 */
            {8'h00}, /* 0x0af6 */
            {8'h00}, /* 0x0af5 */
            {8'h00}, /* 0x0af4 */
            {8'h00}, /* 0x0af3 */
            {8'h00}, /* 0x0af2 */
            {8'h00}, /* 0x0af1 */
            {8'h00}, /* 0x0af0 */
            {8'h00}, /* 0x0aef */
            {8'h00}, /* 0x0aee */
            {8'h00}, /* 0x0aed */
            {8'h00}, /* 0x0aec */
            {8'h00}, /* 0x0aeb */
            {8'h00}, /* 0x0aea */
            {8'h00}, /* 0x0ae9 */
            {8'h00}, /* 0x0ae8 */
            {8'h00}, /* 0x0ae7 */
            {8'h00}, /* 0x0ae6 */
            {8'h00}, /* 0x0ae5 */
            {8'h00}, /* 0x0ae4 */
            {8'h00}, /* 0x0ae3 */
            {8'h00}, /* 0x0ae2 */
            {8'h00}, /* 0x0ae1 */
            {8'h00}, /* 0x0ae0 */
            {8'h00}, /* 0x0adf */
            {8'h00}, /* 0x0ade */
            {8'h00}, /* 0x0add */
            {8'h00}, /* 0x0adc */
            {8'h00}, /* 0x0adb */
            {8'h00}, /* 0x0ada */
            {8'h00}, /* 0x0ad9 */
            {8'h00}, /* 0x0ad8 */
            {8'h00}, /* 0x0ad7 */
            {8'h00}, /* 0x0ad6 */
            {8'h00}, /* 0x0ad5 */
            {8'h00}, /* 0x0ad4 */
            {8'h00}, /* 0x0ad3 */
            {8'h00}, /* 0x0ad2 */
            {8'h00}, /* 0x0ad1 */
            {8'h00}, /* 0x0ad0 */
            {8'h00}, /* 0x0acf */
            {8'h00}, /* 0x0ace */
            {8'h00}, /* 0x0acd */
            {8'h00}, /* 0x0acc */
            {8'h00}, /* 0x0acb */
            {8'h00}, /* 0x0aca */
            {8'h00}, /* 0x0ac9 */
            {8'h00}, /* 0x0ac8 */
            {8'h00}, /* 0x0ac7 */
            {8'h00}, /* 0x0ac6 */
            {8'h00}, /* 0x0ac5 */
            {8'h00}, /* 0x0ac4 */
            {8'h00}, /* 0x0ac3 */
            {8'h00}, /* 0x0ac2 */
            {8'h00}, /* 0x0ac1 */
            {8'h00}, /* 0x0ac0 */
            {8'h00}, /* 0x0abf */
            {8'h00}, /* 0x0abe */
            {8'h00}, /* 0x0abd */
            {8'h00}, /* 0x0abc */
            {8'h00}, /* 0x0abb */
            {8'h00}, /* 0x0aba */
            {8'h00}, /* 0x0ab9 */
            {8'h00}, /* 0x0ab8 */
            {8'h00}, /* 0x0ab7 */
            {8'h00}, /* 0x0ab6 */
            {8'h00}, /* 0x0ab5 */
            {8'h00}, /* 0x0ab4 */
            {8'h00}, /* 0x0ab3 */
            {8'h00}, /* 0x0ab2 */
            {8'h00}, /* 0x0ab1 */
            {8'h00}, /* 0x0ab0 */
            {8'h00}, /* 0x0aaf */
            {8'h00}, /* 0x0aae */
            {8'h00}, /* 0x0aad */
            {8'h00}, /* 0x0aac */
            {8'h00}, /* 0x0aab */
            {8'h00}, /* 0x0aaa */
            {8'h00}, /* 0x0aa9 */
            {8'h00}, /* 0x0aa8 */
            {8'h00}, /* 0x0aa7 */
            {8'h00}, /* 0x0aa6 */
            {8'h00}, /* 0x0aa5 */
            {8'h00}, /* 0x0aa4 */
            {8'h00}, /* 0x0aa3 */
            {8'h00}, /* 0x0aa2 */
            {8'h00}, /* 0x0aa1 */
            {8'h00}, /* 0x0aa0 */
            {8'h00}, /* 0x0a9f */
            {8'h00}, /* 0x0a9e */
            {8'h00}, /* 0x0a9d */
            {8'h00}, /* 0x0a9c */
            {8'h00}, /* 0x0a9b */
            {8'h00}, /* 0x0a9a */
            {8'h00}, /* 0x0a99 */
            {8'h00}, /* 0x0a98 */
            {8'h00}, /* 0x0a97 */
            {8'h00}, /* 0x0a96 */
            {8'h00}, /* 0x0a95 */
            {8'h00}, /* 0x0a94 */
            {8'h00}, /* 0x0a93 */
            {8'h00}, /* 0x0a92 */
            {8'h00}, /* 0x0a91 */
            {8'h00}, /* 0x0a90 */
            {8'h00}, /* 0x0a8f */
            {8'h00}, /* 0x0a8e */
            {8'h00}, /* 0x0a8d */
            {8'h00}, /* 0x0a8c */
            {8'h00}, /* 0x0a8b */
            {8'h00}, /* 0x0a8a */
            {8'h00}, /* 0x0a89 */
            {8'h00}, /* 0x0a88 */
            {8'h00}, /* 0x0a87 */
            {8'h00}, /* 0x0a86 */
            {8'h00}, /* 0x0a85 */
            {8'h00}, /* 0x0a84 */
            {8'h00}, /* 0x0a83 */
            {8'h00}, /* 0x0a82 */
            {8'h00}, /* 0x0a81 */
            {8'h00}, /* 0x0a80 */
            {8'h00}, /* 0x0a7f */
            {8'h00}, /* 0x0a7e */
            {8'h00}, /* 0x0a7d */
            {8'h00}, /* 0x0a7c */
            {8'h00}, /* 0x0a7b */
            {8'h00}, /* 0x0a7a */
            {8'h00}, /* 0x0a79 */
            {8'h00}, /* 0x0a78 */
            {8'h00}, /* 0x0a77 */
            {8'h00}, /* 0x0a76 */
            {8'h00}, /* 0x0a75 */
            {8'h00}, /* 0x0a74 */
            {8'h00}, /* 0x0a73 */
            {8'h00}, /* 0x0a72 */
            {8'h00}, /* 0x0a71 */
            {8'h00}, /* 0x0a70 */
            {8'h00}, /* 0x0a6f */
            {8'h00}, /* 0x0a6e */
            {8'h00}, /* 0x0a6d */
            {8'h00}, /* 0x0a6c */
            {8'h00}, /* 0x0a6b */
            {8'h00}, /* 0x0a6a */
            {8'h00}, /* 0x0a69 */
            {8'h00}, /* 0x0a68 */
            {8'h00}, /* 0x0a67 */
            {8'h00}, /* 0x0a66 */
            {8'h00}, /* 0x0a65 */
            {8'h00}, /* 0x0a64 */
            {8'h00}, /* 0x0a63 */
            {8'h00}, /* 0x0a62 */
            {8'h00}, /* 0x0a61 */
            {8'h00}, /* 0x0a60 */
            {8'h00}, /* 0x0a5f */
            {8'h00}, /* 0x0a5e */
            {8'h00}, /* 0x0a5d */
            {8'h00}, /* 0x0a5c */
            {8'h00}, /* 0x0a5b */
            {8'h00}, /* 0x0a5a */
            {8'h00}, /* 0x0a59 */
            {8'h00}, /* 0x0a58 */
            {8'h00}, /* 0x0a57 */
            {8'h00}, /* 0x0a56 */
            {8'h00}, /* 0x0a55 */
            {8'h00}, /* 0x0a54 */
            {8'h00}, /* 0x0a53 */
            {8'h00}, /* 0x0a52 */
            {8'h00}, /* 0x0a51 */
            {8'h00}, /* 0x0a50 */
            {8'h00}, /* 0x0a4f */
            {8'h00}, /* 0x0a4e */
            {8'h00}, /* 0x0a4d */
            {8'h00}, /* 0x0a4c */
            {8'h00}, /* 0x0a4b */
            {8'h00}, /* 0x0a4a */
            {8'h00}, /* 0x0a49 */
            {8'h00}, /* 0x0a48 */
            {8'h00}, /* 0x0a47 */
            {8'h00}, /* 0x0a46 */
            {8'h00}, /* 0x0a45 */
            {8'h00}, /* 0x0a44 */
            {8'h00}, /* 0x0a43 */
            {8'h00}, /* 0x0a42 */
            {8'h00}, /* 0x0a41 */
            {8'h00}, /* 0x0a40 */
            {8'h00}, /* 0x0a3f */
            {8'h00}, /* 0x0a3e */
            {8'h00}, /* 0x0a3d */
            {8'h00}, /* 0x0a3c */
            {8'h00}, /* 0x0a3b */
            {8'h00}, /* 0x0a3a */
            {8'h00}, /* 0x0a39 */
            {8'h00}, /* 0x0a38 */
            {8'h00}, /* 0x0a37 */
            {8'h00}, /* 0x0a36 */
            {8'h00}, /* 0x0a35 */
            {8'h00}, /* 0x0a34 */
            {8'h00}, /* 0x0a33 */
            {8'h00}, /* 0x0a32 */
            {8'h00}, /* 0x0a31 */
            {8'h00}, /* 0x0a30 */
            {8'h00}, /* 0x0a2f */
            {8'h00}, /* 0x0a2e */
            {8'h00}, /* 0x0a2d */
            {8'h00}, /* 0x0a2c */
            {8'h00}, /* 0x0a2b */
            {8'h00}, /* 0x0a2a */
            {8'h00}, /* 0x0a29 */
            {8'h00}, /* 0x0a28 */
            {8'h00}, /* 0x0a27 */
            {8'h00}, /* 0x0a26 */
            {8'h00}, /* 0x0a25 */
            {8'h00}, /* 0x0a24 */
            {8'h00}, /* 0x0a23 */
            {8'h00}, /* 0x0a22 */
            {8'h00}, /* 0x0a21 */
            {8'h00}, /* 0x0a20 */
            {8'h00}, /* 0x0a1f */
            {8'h00}, /* 0x0a1e */
            {8'h00}, /* 0x0a1d */
            {8'h00}, /* 0x0a1c */
            {8'h00}, /* 0x0a1b */
            {8'h00}, /* 0x0a1a */
            {8'h00}, /* 0x0a19 */
            {8'h00}, /* 0x0a18 */
            {8'h00}, /* 0x0a17 */
            {8'h00}, /* 0x0a16 */
            {8'h00}, /* 0x0a15 */
            {8'h00}, /* 0x0a14 */
            {8'h00}, /* 0x0a13 */
            {8'h00}, /* 0x0a12 */
            {8'h00}, /* 0x0a11 */
            {8'h00}, /* 0x0a10 */
            {8'h00}, /* 0x0a0f */
            {8'h00}, /* 0x0a0e */
            {8'h00}, /* 0x0a0d */
            {8'h00}, /* 0x0a0c */
            {8'h00}, /* 0x0a0b */
            {8'h00}, /* 0x0a0a */
            {8'h00}, /* 0x0a09 */
            {8'h00}, /* 0x0a08 */
            {8'h00}, /* 0x0a07 */
            {8'h00}, /* 0x0a06 */
            {8'h00}, /* 0x0a05 */
            {8'h00}, /* 0x0a04 */
            {8'h00}, /* 0x0a03 */
            {8'h00}, /* 0x0a02 */
            {8'h00}, /* 0x0a01 */
            {8'h00}, /* 0x0a00 */
            {8'h00}, /* 0x09ff */
            {8'h00}, /* 0x09fe */
            {8'h00}, /* 0x09fd */
            {8'h00}, /* 0x09fc */
            {8'h00}, /* 0x09fb */
            {8'h00}, /* 0x09fa */
            {8'h00}, /* 0x09f9 */
            {8'h00}, /* 0x09f8 */
            {8'h00}, /* 0x09f7 */
            {8'h00}, /* 0x09f6 */
            {8'h00}, /* 0x09f5 */
            {8'h00}, /* 0x09f4 */
            {8'h00}, /* 0x09f3 */
            {8'h00}, /* 0x09f2 */
            {8'h00}, /* 0x09f1 */
            {8'h00}, /* 0x09f0 */
            {8'h00}, /* 0x09ef */
            {8'h00}, /* 0x09ee */
            {8'h00}, /* 0x09ed */
            {8'h00}, /* 0x09ec */
            {8'h00}, /* 0x09eb */
            {8'h00}, /* 0x09ea */
            {8'h00}, /* 0x09e9 */
            {8'h00}, /* 0x09e8 */
            {8'h00}, /* 0x09e7 */
            {8'h00}, /* 0x09e6 */
            {8'h00}, /* 0x09e5 */
            {8'h00}, /* 0x09e4 */
            {8'h00}, /* 0x09e3 */
            {8'h00}, /* 0x09e2 */
            {8'h00}, /* 0x09e1 */
            {8'h00}, /* 0x09e0 */
            {8'h00}, /* 0x09df */
            {8'h00}, /* 0x09de */
            {8'h00}, /* 0x09dd */
            {8'h00}, /* 0x09dc */
            {8'h00}, /* 0x09db */
            {8'h00}, /* 0x09da */
            {8'h00}, /* 0x09d9 */
            {8'h00}, /* 0x09d8 */
            {8'h00}, /* 0x09d7 */
            {8'h00}, /* 0x09d6 */
            {8'h00}, /* 0x09d5 */
            {8'h00}, /* 0x09d4 */
            {8'h00}, /* 0x09d3 */
            {8'h00}, /* 0x09d2 */
            {8'h00}, /* 0x09d1 */
            {8'h00}, /* 0x09d0 */
            {8'h00}, /* 0x09cf */
            {8'h00}, /* 0x09ce */
            {8'h00}, /* 0x09cd */
            {8'h00}, /* 0x09cc */
            {8'h00}, /* 0x09cb */
            {8'h00}, /* 0x09ca */
            {8'h00}, /* 0x09c9 */
            {8'h00}, /* 0x09c8 */
            {8'h00}, /* 0x09c7 */
            {8'h00}, /* 0x09c6 */
            {8'h00}, /* 0x09c5 */
            {8'h00}, /* 0x09c4 */
            {8'h00}, /* 0x09c3 */
            {8'h00}, /* 0x09c2 */
            {8'h00}, /* 0x09c1 */
            {8'h00}, /* 0x09c0 */
            {8'h00}, /* 0x09bf */
            {8'h00}, /* 0x09be */
            {8'h00}, /* 0x09bd */
            {8'h00}, /* 0x09bc */
            {8'h00}, /* 0x09bb */
            {8'h00}, /* 0x09ba */
            {8'h00}, /* 0x09b9 */
            {8'h00}, /* 0x09b8 */
            {8'h00}, /* 0x09b7 */
            {8'h00}, /* 0x09b6 */
            {8'h00}, /* 0x09b5 */
            {8'h00}, /* 0x09b4 */
            {8'h00}, /* 0x09b3 */
            {8'h00}, /* 0x09b2 */
            {8'h00}, /* 0x09b1 */
            {8'h00}, /* 0x09b0 */
            {8'h00}, /* 0x09af */
            {8'h00}, /* 0x09ae */
            {8'h00}, /* 0x09ad */
            {8'h00}, /* 0x09ac */
            {8'h00}, /* 0x09ab */
            {8'h00}, /* 0x09aa */
            {8'h00}, /* 0x09a9 */
            {8'h00}, /* 0x09a8 */
            {8'h00}, /* 0x09a7 */
            {8'h00}, /* 0x09a6 */
            {8'h00}, /* 0x09a5 */
            {8'h00}, /* 0x09a4 */
            {8'h00}, /* 0x09a3 */
            {8'h00}, /* 0x09a2 */
            {8'h00}, /* 0x09a1 */
            {8'h00}, /* 0x09a0 */
            {8'h00}, /* 0x099f */
            {8'h00}, /* 0x099e */
            {8'h00}, /* 0x099d */
            {8'h00}, /* 0x099c */
            {8'h00}, /* 0x099b */
            {8'h00}, /* 0x099a */
            {8'h00}, /* 0x0999 */
            {8'h00}, /* 0x0998 */
            {8'h00}, /* 0x0997 */
            {8'h00}, /* 0x0996 */
            {8'h00}, /* 0x0995 */
            {8'h00}, /* 0x0994 */
            {8'h00}, /* 0x0993 */
            {8'h00}, /* 0x0992 */
            {8'h00}, /* 0x0991 */
            {8'h00}, /* 0x0990 */
            {8'h00}, /* 0x098f */
            {8'h00}, /* 0x098e */
            {8'h00}, /* 0x098d */
            {8'h00}, /* 0x098c */
            {8'h00}, /* 0x098b */
            {8'h00}, /* 0x098a */
            {8'h00}, /* 0x0989 */
            {8'h00}, /* 0x0988 */
            {8'h00}, /* 0x0987 */
            {8'h00}, /* 0x0986 */
            {8'h00}, /* 0x0985 */
            {8'h00}, /* 0x0984 */
            {8'h00}, /* 0x0983 */
            {8'h00}, /* 0x0982 */
            {8'h00}, /* 0x0981 */
            {8'h00}, /* 0x0980 */
            {8'h00}, /* 0x097f */
            {8'h00}, /* 0x097e */
            {8'h00}, /* 0x097d */
            {8'h00}, /* 0x097c */
            {8'h00}, /* 0x097b */
            {8'h00}, /* 0x097a */
            {8'h00}, /* 0x0979 */
            {8'h00}, /* 0x0978 */
            {8'h00}, /* 0x0977 */
            {8'h00}, /* 0x0976 */
            {8'h00}, /* 0x0975 */
            {8'h00}, /* 0x0974 */
            {8'h00}, /* 0x0973 */
            {8'h00}, /* 0x0972 */
            {8'h00}, /* 0x0971 */
            {8'h00}, /* 0x0970 */
            {8'h00}, /* 0x096f */
            {8'h00}, /* 0x096e */
            {8'h00}, /* 0x096d */
            {8'h00}, /* 0x096c */
            {8'h00}, /* 0x096b */
            {8'h00}, /* 0x096a */
            {8'h00}, /* 0x0969 */
            {8'h00}, /* 0x0968 */
            {8'h00}, /* 0x0967 */
            {8'h00}, /* 0x0966 */
            {8'h00}, /* 0x0965 */
            {8'h00}, /* 0x0964 */
            {8'h00}, /* 0x0963 */
            {8'h00}, /* 0x0962 */
            {8'h00}, /* 0x0961 */
            {8'h00}, /* 0x0960 */
            {8'h00}, /* 0x095f */
            {8'h00}, /* 0x095e */
            {8'h00}, /* 0x095d */
            {8'h00}, /* 0x095c */
            {8'h00}, /* 0x095b */
            {8'h00}, /* 0x095a */
            {8'h00}, /* 0x0959 */
            {8'h00}, /* 0x0958 */
            {8'h00}, /* 0x0957 */
            {8'h00}, /* 0x0956 */
            {8'h00}, /* 0x0955 */
            {8'h00}, /* 0x0954 */
            {8'h00}, /* 0x0953 */
            {8'h00}, /* 0x0952 */
            {8'h00}, /* 0x0951 */
            {8'h00}, /* 0x0950 */
            {8'h00}, /* 0x094f */
            {8'h00}, /* 0x094e */
            {8'h00}, /* 0x094d */
            {8'h00}, /* 0x094c */
            {8'h00}, /* 0x094b */
            {8'h00}, /* 0x094a */
            {8'h00}, /* 0x0949 */
            {8'h00}, /* 0x0948 */
            {8'h00}, /* 0x0947 */
            {8'h00}, /* 0x0946 */
            {8'h00}, /* 0x0945 */
            {8'h00}, /* 0x0944 */
            {8'h00}, /* 0x0943 */
            {8'h00}, /* 0x0942 */
            {8'h00}, /* 0x0941 */
            {8'h00}, /* 0x0940 */
            {8'h00}, /* 0x093f */
            {8'h00}, /* 0x093e */
            {8'h00}, /* 0x093d */
            {8'h00}, /* 0x093c */
            {8'h00}, /* 0x093b */
            {8'h00}, /* 0x093a */
            {8'h00}, /* 0x0939 */
            {8'h00}, /* 0x0938 */
            {8'h00}, /* 0x0937 */
            {8'h00}, /* 0x0936 */
            {8'h00}, /* 0x0935 */
            {8'h00}, /* 0x0934 */
            {8'h00}, /* 0x0933 */
            {8'h00}, /* 0x0932 */
            {8'h00}, /* 0x0931 */
            {8'h00}, /* 0x0930 */
            {8'h00}, /* 0x092f */
            {8'h00}, /* 0x092e */
            {8'h00}, /* 0x092d */
            {8'h00}, /* 0x092c */
            {8'h00}, /* 0x092b */
            {8'h00}, /* 0x092a */
            {8'h00}, /* 0x0929 */
            {8'h00}, /* 0x0928 */
            {8'h00}, /* 0x0927 */
            {8'h00}, /* 0x0926 */
            {8'h00}, /* 0x0925 */
            {8'h00}, /* 0x0924 */
            {8'h00}, /* 0x0923 */
            {8'h00}, /* 0x0922 */
            {8'h00}, /* 0x0921 */
            {8'h00}, /* 0x0920 */
            {8'h00}, /* 0x091f */
            {8'h00}, /* 0x091e */
            {8'h00}, /* 0x091d */
            {8'h00}, /* 0x091c */
            {8'h00}, /* 0x091b */
            {8'h00}, /* 0x091a */
            {8'h00}, /* 0x0919 */
            {8'h00}, /* 0x0918 */
            {8'h00}, /* 0x0917 */
            {8'h00}, /* 0x0916 */
            {8'h00}, /* 0x0915 */
            {8'h00}, /* 0x0914 */
            {8'h00}, /* 0x0913 */
            {8'h00}, /* 0x0912 */
            {8'h00}, /* 0x0911 */
            {8'h00}, /* 0x0910 */
            {8'h00}, /* 0x090f */
            {8'h00}, /* 0x090e */
            {8'h00}, /* 0x090d */
            {8'h00}, /* 0x090c */
            {8'h00}, /* 0x090b */
            {8'h00}, /* 0x090a */
            {8'h00}, /* 0x0909 */
            {8'h00}, /* 0x0908 */
            {8'h00}, /* 0x0907 */
            {8'h00}, /* 0x0906 */
            {8'h00}, /* 0x0905 */
            {8'h00}, /* 0x0904 */
            {8'h00}, /* 0x0903 */
            {8'h00}, /* 0x0902 */
            {8'h00}, /* 0x0901 */
            {8'h00}, /* 0x0900 */
            {8'h00}, /* 0x08ff */
            {8'h00}, /* 0x08fe */
            {8'h00}, /* 0x08fd */
            {8'h00}, /* 0x08fc */
            {8'h00}, /* 0x08fb */
            {8'h00}, /* 0x08fa */
            {8'h00}, /* 0x08f9 */
            {8'h00}, /* 0x08f8 */
            {8'h00}, /* 0x08f7 */
            {8'h00}, /* 0x08f6 */
            {8'h00}, /* 0x08f5 */
            {8'h00}, /* 0x08f4 */
            {8'h00}, /* 0x08f3 */
            {8'h00}, /* 0x08f2 */
            {8'h00}, /* 0x08f1 */
            {8'h00}, /* 0x08f0 */
            {8'h00}, /* 0x08ef */
            {8'h00}, /* 0x08ee */
            {8'h00}, /* 0x08ed */
            {8'h00}, /* 0x08ec */
            {8'h00}, /* 0x08eb */
            {8'h00}, /* 0x08ea */
            {8'h00}, /* 0x08e9 */
            {8'h00}, /* 0x08e8 */
            {8'h00}, /* 0x08e7 */
            {8'h00}, /* 0x08e6 */
            {8'h00}, /* 0x08e5 */
            {8'h00}, /* 0x08e4 */
            {8'h00}, /* 0x08e3 */
            {8'h00}, /* 0x08e2 */
            {8'h00}, /* 0x08e1 */
            {8'h00}, /* 0x08e0 */
            {8'h00}, /* 0x08df */
            {8'h00}, /* 0x08de */
            {8'h00}, /* 0x08dd */
            {8'h00}, /* 0x08dc */
            {8'h00}, /* 0x08db */
            {8'h00}, /* 0x08da */
            {8'h00}, /* 0x08d9 */
            {8'h00}, /* 0x08d8 */
            {8'h00}, /* 0x08d7 */
            {8'h00}, /* 0x08d6 */
            {8'h00}, /* 0x08d5 */
            {8'h00}, /* 0x08d4 */
            {8'h00}, /* 0x08d3 */
            {8'h00}, /* 0x08d2 */
            {8'h00}, /* 0x08d1 */
            {8'h00}, /* 0x08d0 */
            {8'h00}, /* 0x08cf */
            {8'h00}, /* 0x08ce */
            {8'h00}, /* 0x08cd */
            {8'h00}, /* 0x08cc */
            {8'h00}, /* 0x08cb */
            {8'h00}, /* 0x08ca */
            {8'h00}, /* 0x08c9 */
            {8'h00}, /* 0x08c8 */
            {8'h00}, /* 0x08c7 */
            {8'h00}, /* 0x08c6 */
            {8'h00}, /* 0x08c5 */
            {8'h00}, /* 0x08c4 */
            {8'h00}, /* 0x08c3 */
            {8'h00}, /* 0x08c2 */
            {8'h00}, /* 0x08c1 */
            {8'h00}, /* 0x08c0 */
            {8'h00}, /* 0x08bf */
            {8'h00}, /* 0x08be */
            {8'h00}, /* 0x08bd */
            {8'h00}, /* 0x08bc */
            {8'h00}, /* 0x08bb */
            {8'h00}, /* 0x08ba */
            {8'h00}, /* 0x08b9 */
            {8'h00}, /* 0x08b8 */
            {8'h00}, /* 0x08b7 */
            {8'h00}, /* 0x08b6 */
            {8'h00}, /* 0x08b5 */
            {8'h00}, /* 0x08b4 */
            {8'h00}, /* 0x08b3 */
            {8'h00}, /* 0x08b2 */
            {8'h00}, /* 0x08b1 */
            {8'h00}, /* 0x08b0 */
            {8'h00}, /* 0x08af */
            {8'h00}, /* 0x08ae */
            {8'h00}, /* 0x08ad */
            {8'h00}, /* 0x08ac */
            {8'h00}, /* 0x08ab */
            {8'h00}, /* 0x08aa */
            {8'h00}, /* 0x08a9 */
            {8'h00}, /* 0x08a8 */
            {8'h00}, /* 0x08a7 */
            {8'h00}, /* 0x08a6 */
            {8'h00}, /* 0x08a5 */
            {8'h00}, /* 0x08a4 */
            {8'h00}, /* 0x08a3 */
            {8'h00}, /* 0x08a2 */
            {8'h00}, /* 0x08a1 */
            {8'h00}, /* 0x08a0 */
            {8'h00}, /* 0x089f */
            {8'h00}, /* 0x089e */
            {8'h00}, /* 0x089d */
            {8'h00}, /* 0x089c */
            {8'h00}, /* 0x089b */
            {8'h00}, /* 0x089a */
            {8'h00}, /* 0x0899 */
            {8'h00}, /* 0x0898 */
            {8'h00}, /* 0x0897 */
            {8'h00}, /* 0x0896 */
            {8'h00}, /* 0x0895 */
            {8'h00}, /* 0x0894 */
            {8'h00}, /* 0x0893 */
            {8'h00}, /* 0x0892 */
            {8'h00}, /* 0x0891 */
            {8'h00}, /* 0x0890 */
            {8'h00}, /* 0x088f */
            {8'h00}, /* 0x088e */
            {8'h00}, /* 0x088d */
            {8'h00}, /* 0x088c */
            {8'h00}, /* 0x088b */
            {8'h00}, /* 0x088a */
            {8'h00}, /* 0x0889 */
            {8'h00}, /* 0x0888 */
            {8'h00}, /* 0x0887 */
            {8'h00}, /* 0x0886 */
            {8'h00}, /* 0x0885 */
            {8'h00}, /* 0x0884 */
            {8'h00}, /* 0x0883 */
            {8'h00}, /* 0x0882 */
            {8'h00}, /* 0x0881 */
            {8'h00}, /* 0x0880 */
            {8'h00}, /* 0x087f */
            {8'h00}, /* 0x087e */
            {8'h00}, /* 0x087d */
            {8'h00}, /* 0x087c */
            {8'h00}, /* 0x087b */
            {8'h00}, /* 0x087a */
            {8'h00}, /* 0x0879 */
            {8'h00}, /* 0x0878 */
            {8'h00}, /* 0x0877 */
            {8'h00}, /* 0x0876 */
            {8'h00}, /* 0x0875 */
            {8'h00}, /* 0x0874 */
            {8'h00}, /* 0x0873 */
            {8'h00}, /* 0x0872 */
            {8'h00}, /* 0x0871 */
            {8'h00}, /* 0x0870 */
            {8'h00}, /* 0x086f */
            {8'h00}, /* 0x086e */
            {8'h00}, /* 0x086d */
            {8'h00}, /* 0x086c */
            {8'h00}, /* 0x086b */
            {8'h00}, /* 0x086a */
            {8'h00}, /* 0x0869 */
            {8'h00}, /* 0x0868 */
            {8'h00}, /* 0x0867 */
            {8'h00}, /* 0x0866 */
            {8'h00}, /* 0x0865 */
            {8'h00}, /* 0x0864 */
            {8'h00}, /* 0x0863 */
            {8'h00}, /* 0x0862 */
            {8'h00}, /* 0x0861 */
            {8'h00}, /* 0x0860 */
            {8'h00}, /* 0x085f */
            {8'h00}, /* 0x085e */
            {8'h00}, /* 0x085d */
            {8'h00}, /* 0x085c */
            {8'h00}, /* 0x085b */
            {8'h00}, /* 0x085a */
            {8'h00}, /* 0x0859 */
            {8'h00}, /* 0x0858 */
            {8'h00}, /* 0x0857 */
            {8'h00}, /* 0x0856 */
            {8'h00}, /* 0x0855 */
            {8'h00}, /* 0x0854 */
            {8'h00}, /* 0x0853 */
            {8'h00}, /* 0x0852 */
            {8'h00}, /* 0x0851 */
            {8'h00}, /* 0x0850 */
            {8'h00}, /* 0x084f */
            {8'h00}, /* 0x084e */
            {8'h00}, /* 0x084d */
            {8'h00}, /* 0x084c */
            {8'h00}, /* 0x084b */
            {8'h00}, /* 0x084a */
            {8'h00}, /* 0x0849 */
            {8'h00}, /* 0x0848 */
            {8'h00}, /* 0x0847 */
            {8'h00}, /* 0x0846 */
            {8'h00}, /* 0x0845 */
            {8'h00}, /* 0x0844 */
            {8'h00}, /* 0x0843 */
            {8'h00}, /* 0x0842 */
            {8'h00}, /* 0x0841 */
            {8'h00}, /* 0x0840 */
            {8'h00}, /* 0x083f */
            {8'h00}, /* 0x083e */
            {8'h00}, /* 0x083d */
            {8'h00}, /* 0x083c */
            {8'h00}, /* 0x083b */
            {8'h00}, /* 0x083a */
            {8'h00}, /* 0x0839 */
            {8'h00}, /* 0x0838 */
            {8'h00}, /* 0x0837 */
            {8'h00}, /* 0x0836 */
            {8'h00}, /* 0x0835 */
            {8'h00}, /* 0x0834 */
            {8'h00}, /* 0x0833 */
            {8'h00}, /* 0x0832 */
            {8'h00}, /* 0x0831 */
            {8'h00}, /* 0x0830 */
            {8'h00}, /* 0x082f */
            {8'h00}, /* 0x082e */
            {8'h00}, /* 0x082d */
            {8'h00}, /* 0x082c */
            {8'h00}, /* 0x082b */
            {8'h00}, /* 0x082a */
            {8'h00}, /* 0x0829 */
            {8'h00}, /* 0x0828 */
            {8'h00}, /* 0x0827 */
            {8'h00}, /* 0x0826 */
            {8'h00}, /* 0x0825 */
            {8'h00}, /* 0x0824 */
            {8'h00}, /* 0x0823 */
            {8'h00}, /* 0x0822 */
            {8'h00}, /* 0x0821 */
            {8'h00}, /* 0x0820 */
            {8'h00}, /* 0x081f */
            {8'h00}, /* 0x081e */
            {8'h00}, /* 0x081d */
            {8'h00}, /* 0x081c */
            {8'h00}, /* 0x081b */
            {8'h00}, /* 0x081a */
            {8'h00}, /* 0x0819 */
            {8'h00}, /* 0x0818 */
            {8'h00}, /* 0x0817 */
            {8'h00}, /* 0x0816 */
            {8'h00}, /* 0x0815 */
            {8'h00}, /* 0x0814 */
            {8'h00}, /* 0x0813 */
            {8'h00}, /* 0x0812 */
            {8'h00}, /* 0x0811 */
            {8'h00}, /* 0x0810 */
            {8'h00}, /* 0x080f */
            {8'h00}, /* 0x080e */
            {8'h00}, /* 0x080d */
            {8'h00}, /* 0x080c */
            {8'h00}, /* 0x080b */
            {8'h00}, /* 0x080a */
            {8'h00}, /* 0x0809 */
            {8'h00}, /* 0x0808 */
            {8'h00}, /* 0x0807 */
            {8'h00}, /* 0x0806 */
            {8'h00}, /* 0x0805 */
            {8'h00}, /* 0x0804 */
            {8'h00}, /* 0x0803 */
            {8'h00}, /* 0x0802 */
            {8'h00}, /* 0x0801 */
            {8'h00}, /* 0x0800 */
            {8'h00}, /* 0x07ff */
            {8'h00}, /* 0x07fe */
            {8'h00}, /* 0x07fd */
            {8'h00}, /* 0x07fc */
            {8'h00}, /* 0x07fb */
            {8'h00}, /* 0x07fa */
            {8'h00}, /* 0x07f9 */
            {8'h00}, /* 0x07f8 */
            {8'h00}, /* 0x07f7 */
            {8'h00}, /* 0x07f6 */
            {8'h00}, /* 0x07f5 */
            {8'h00}, /* 0x07f4 */
            {8'h00}, /* 0x07f3 */
            {8'h00}, /* 0x07f2 */
            {8'h00}, /* 0x07f1 */
            {8'h00}, /* 0x07f0 */
            {8'h00}, /* 0x07ef */
            {8'h00}, /* 0x07ee */
            {8'h00}, /* 0x07ed */
            {8'h00}, /* 0x07ec */
            {8'h00}, /* 0x07eb */
            {8'h00}, /* 0x07ea */
            {8'h00}, /* 0x07e9 */
            {8'h00}, /* 0x07e8 */
            {8'h00}, /* 0x07e7 */
            {8'h00}, /* 0x07e6 */
            {8'h00}, /* 0x07e5 */
            {8'h00}, /* 0x07e4 */
            {8'h00}, /* 0x07e3 */
            {8'h00}, /* 0x07e2 */
            {8'h00}, /* 0x07e1 */
            {8'h00}, /* 0x07e0 */
            {8'h00}, /* 0x07df */
            {8'h00}, /* 0x07de */
            {8'h00}, /* 0x07dd */
            {8'h00}, /* 0x07dc */
            {8'h00}, /* 0x07db */
            {8'h00}, /* 0x07da */
            {8'h00}, /* 0x07d9 */
            {8'h00}, /* 0x07d8 */
            {8'h00}, /* 0x07d7 */
            {8'h00}, /* 0x07d6 */
            {8'h00}, /* 0x07d5 */
            {8'h00}, /* 0x07d4 */
            {8'h00}, /* 0x07d3 */
            {8'h00}, /* 0x07d2 */
            {8'h00}, /* 0x07d1 */
            {8'h00}, /* 0x07d0 */
            {8'h00}, /* 0x07cf */
            {8'h00}, /* 0x07ce */
            {8'h00}, /* 0x07cd */
            {8'h00}, /* 0x07cc */
            {8'h00}, /* 0x07cb */
            {8'h00}, /* 0x07ca */
            {8'h00}, /* 0x07c9 */
            {8'h00}, /* 0x07c8 */
            {8'h00}, /* 0x07c7 */
            {8'h00}, /* 0x07c6 */
            {8'h00}, /* 0x07c5 */
            {8'h00}, /* 0x07c4 */
            {8'h00}, /* 0x07c3 */
            {8'h00}, /* 0x07c2 */
            {8'h00}, /* 0x07c1 */
            {8'h00}, /* 0x07c0 */
            {8'h00}, /* 0x07bf */
            {8'h00}, /* 0x07be */
            {8'h00}, /* 0x07bd */
            {8'h00}, /* 0x07bc */
            {8'h00}, /* 0x07bb */
            {8'h00}, /* 0x07ba */
            {8'h00}, /* 0x07b9 */
            {8'h00}, /* 0x07b8 */
            {8'h00}, /* 0x07b7 */
            {8'h00}, /* 0x07b6 */
            {8'h00}, /* 0x07b5 */
            {8'h00}, /* 0x07b4 */
            {8'h00}, /* 0x07b3 */
            {8'h00}, /* 0x07b2 */
            {8'h00}, /* 0x07b1 */
            {8'h00}, /* 0x07b0 */
            {8'h00}, /* 0x07af */
            {8'h00}, /* 0x07ae */
            {8'h00}, /* 0x07ad */
            {8'h00}, /* 0x07ac */
            {8'h00}, /* 0x07ab */
            {8'h00}, /* 0x07aa */
            {8'h00}, /* 0x07a9 */
            {8'h00}, /* 0x07a8 */
            {8'h00}, /* 0x07a7 */
            {8'h00}, /* 0x07a6 */
            {8'h00}, /* 0x07a5 */
            {8'h00}, /* 0x07a4 */
            {8'h00}, /* 0x07a3 */
            {8'h00}, /* 0x07a2 */
            {8'h00}, /* 0x07a1 */
            {8'h00}, /* 0x07a0 */
            {8'h00}, /* 0x079f */
            {8'h00}, /* 0x079e */
            {8'h00}, /* 0x079d */
            {8'h00}, /* 0x079c */
            {8'h00}, /* 0x079b */
            {8'h00}, /* 0x079a */
            {8'h00}, /* 0x0799 */
            {8'h00}, /* 0x0798 */
            {8'h00}, /* 0x0797 */
            {8'h00}, /* 0x0796 */
            {8'h00}, /* 0x0795 */
            {8'h00}, /* 0x0794 */
            {8'h00}, /* 0x0793 */
            {8'h00}, /* 0x0792 */
            {8'h00}, /* 0x0791 */
            {8'h00}, /* 0x0790 */
            {8'h00}, /* 0x078f */
            {8'h00}, /* 0x078e */
            {8'h00}, /* 0x078d */
            {8'h00}, /* 0x078c */
            {8'h00}, /* 0x078b */
            {8'h00}, /* 0x078a */
            {8'h00}, /* 0x0789 */
            {8'h00}, /* 0x0788 */
            {8'h00}, /* 0x0787 */
            {8'h00}, /* 0x0786 */
            {8'h00}, /* 0x0785 */
            {8'h00}, /* 0x0784 */
            {8'h00}, /* 0x0783 */
            {8'h00}, /* 0x0782 */
            {8'h00}, /* 0x0781 */
            {8'h00}, /* 0x0780 */
            {8'h00}, /* 0x077f */
            {8'h00}, /* 0x077e */
            {8'h00}, /* 0x077d */
            {8'h00}, /* 0x077c */
            {8'h00}, /* 0x077b */
            {8'h00}, /* 0x077a */
            {8'h00}, /* 0x0779 */
            {8'h00}, /* 0x0778 */
            {8'h00}, /* 0x0777 */
            {8'h00}, /* 0x0776 */
            {8'h00}, /* 0x0775 */
            {8'h00}, /* 0x0774 */
            {8'h00}, /* 0x0773 */
            {8'h00}, /* 0x0772 */
            {8'h00}, /* 0x0771 */
            {8'h00}, /* 0x0770 */
            {8'h00}, /* 0x076f */
            {8'h00}, /* 0x076e */
            {8'h00}, /* 0x076d */
            {8'h00}, /* 0x076c */
            {8'h00}, /* 0x076b */
            {8'h00}, /* 0x076a */
            {8'h00}, /* 0x0769 */
            {8'h00}, /* 0x0768 */
            {8'h00}, /* 0x0767 */
            {8'h00}, /* 0x0766 */
            {8'h00}, /* 0x0765 */
            {8'h00}, /* 0x0764 */
            {8'h00}, /* 0x0763 */
            {8'h00}, /* 0x0762 */
            {8'h00}, /* 0x0761 */
            {8'h00}, /* 0x0760 */
            {8'h00}, /* 0x075f */
            {8'h00}, /* 0x075e */
            {8'h00}, /* 0x075d */
            {8'h00}, /* 0x075c */
            {8'h00}, /* 0x075b */
            {8'h00}, /* 0x075a */
            {8'h00}, /* 0x0759 */
            {8'h00}, /* 0x0758 */
            {8'h00}, /* 0x0757 */
            {8'h00}, /* 0x0756 */
            {8'h00}, /* 0x0755 */
            {8'h00}, /* 0x0754 */
            {8'h00}, /* 0x0753 */
            {8'h00}, /* 0x0752 */
            {8'h00}, /* 0x0751 */
            {8'h00}, /* 0x0750 */
            {8'h00}, /* 0x074f */
            {8'h00}, /* 0x074e */
            {8'h00}, /* 0x074d */
            {8'h00}, /* 0x074c */
            {8'h00}, /* 0x074b */
            {8'h00}, /* 0x074a */
            {8'h00}, /* 0x0749 */
            {8'h00}, /* 0x0748 */
            {8'h00}, /* 0x0747 */
            {8'h00}, /* 0x0746 */
            {8'h00}, /* 0x0745 */
            {8'h00}, /* 0x0744 */
            {8'h00}, /* 0x0743 */
            {8'h00}, /* 0x0742 */
            {8'h00}, /* 0x0741 */
            {8'h00}, /* 0x0740 */
            {8'h00}, /* 0x073f */
            {8'h00}, /* 0x073e */
            {8'h00}, /* 0x073d */
            {8'h00}, /* 0x073c */
            {8'h00}, /* 0x073b */
            {8'h00}, /* 0x073a */
            {8'h00}, /* 0x0739 */
            {8'h00}, /* 0x0738 */
            {8'h00}, /* 0x0737 */
            {8'h00}, /* 0x0736 */
            {8'h00}, /* 0x0735 */
            {8'h00}, /* 0x0734 */
            {8'h00}, /* 0x0733 */
            {8'h00}, /* 0x0732 */
            {8'h00}, /* 0x0731 */
            {8'h00}, /* 0x0730 */
            {8'h00}, /* 0x072f */
            {8'h00}, /* 0x072e */
            {8'h00}, /* 0x072d */
            {8'h00}, /* 0x072c */
            {8'h00}, /* 0x072b */
            {8'h00}, /* 0x072a */
            {8'h00}, /* 0x0729 */
            {8'h00}, /* 0x0728 */
            {8'h00}, /* 0x0727 */
            {8'h00}, /* 0x0726 */
            {8'h00}, /* 0x0725 */
            {8'h00}, /* 0x0724 */
            {8'h00}, /* 0x0723 */
            {8'h00}, /* 0x0722 */
            {8'h00}, /* 0x0721 */
            {8'h00}, /* 0x0720 */
            {8'h00}, /* 0x071f */
            {8'h00}, /* 0x071e */
            {8'h00}, /* 0x071d */
            {8'h00}, /* 0x071c */
            {8'h00}, /* 0x071b */
            {8'h00}, /* 0x071a */
            {8'h00}, /* 0x0719 */
            {8'h00}, /* 0x0718 */
            {8'h00}, /* 0x0717 */
            {8'h00}, /* 0x0716 */
            {8'h00}, /* 0x0715 */
            {8'h00}, /* 0x0714 */
            {8'h00}, /* 0x0713 */
            {8'h00}, /* 0x0712 */
            {8'h00}, /* 0x0711 */
            {8'h00}, /* 0x0710 */
            {8'h00}, /* 0x070f */
            {8'h00}, /* 0x070e */
            {8'h00}, /* 0x070d */
            {8'h00}, /* 0x070c */
            {8'h00}, /* 0x070b */
            {8'h00}, /* 0x070a */
            {8'h00}, /* 0x0709 */
            {8'h00}, /* 0x0708 */
            {8'h00}, /* 0x0707 */
            {8'h00}, /* 0x0706 */
            {8'h00}, /* 0x0705 */
            {8'h00}, /* 0x0704 */
            {8'h00}, /* 0x0703 */
            {8'h00}, /* 0x0702 */
            {8'h00}, /* 0x0701 */
            {8'h00}, /* 0x0700 */
            {8'h00}, /* 0x06ff */
            {8'h00}, /* 0x06fe */
            {8'h00}, /* 0x06fd */
            {8'h00}, /* 0x06fc */
            {8'h00}, /* 0x06fb */
            {8'h00}, /* 0x06fa */
            {8'h00}, /* 0x06f9 */
            {8'h00}, /* 0x06f8 */
            {8'h00}, /* 0x06f7 */
            {8'h00}, /* 0x06f6 */
            {8'h00}, /* 0x06f5 */
            {8'h00}, /* 0x06f4 */
            {8'h00}, /* 0x06f3 */
            {8'h00}, /* 0x06f2 */
            {8'h00}, /* 0x06f1 */
            {8'h00}, /* 0x06f0 */
            {8'h00}, /* 0x06ef */
            {8'h00}, /* 0x06ee */
            {8'h00}, /* 0x06ed */
            {8'h00}, /* 0x06ec */
            {8'h00}, /* 0x06eb */
            {8'h00}, /* 0x06ea */
            {8'h00}, /* 0x06e9 */
            {8'h00}, /* 0x06e8 */
            {8'h00}, /* 0x06e7 */
            {8'h00}, /* 0x06e6 */
            {8'h00}, /* 0x06e5 */
            {8'h00}, /* 0x06e4 */
            {8'h00}, /* 0x06e3 */
            {8'h00}, /* 0x06e2 */
            {8'h00}, /* 0x06e1 */
            {8'h00}, /* 0x06e0 */
            {8'h00}, /* 0x06df */
            {8'h00}, /* 0x06de */
            {8'h00}, /* 0x06dd */
            {8'h00}, /* 0x06dc */
            {8'h00}, /* 0x06db */
            {8'h00}, /* 0x06da */
            {8'h00}, /* 0x06d9 */
            {8'h00}, /* 0x06d8 */
            {8'h00}, /* 0x06d7 */
            {8'h00}, /* 0x06d6 */
            {8'h00}, /* 0x06d5 */
            {8'h00}, /* 0x06d4 */
            {8'h00}, /* 0x06d3 */
            {8'h00}, /* 0x06d2 */
            {8'h00}, /* 0x06d1 */
            {8'h00}, /* 0x06d0 */
            {8'h00}, /* 0x06cf */
            {8'h00}, /* 0x06ce */
            {8'h00}, /* 0x06cd */
            {8'h00}, /* 0x06cc */
            {8'h00}, /* 0x06cb */
            {8'h00}, /* 0x06ca */
            {8'h00}, /* 0x06c9 */
            {8'h00}, /* 0x06c8 */
            {8'h00}, /* 0x06c7 */
            {8'h00}, /* 0x06c6 */
            {8'h00}, /* 0x06c5 */
            {8'h00}, /* 0x06c4 */
            {8'h00}, /* 0x06c3 */
            {8'h00}, /* 0x06c2 */
            {8'h00}, /* 0x06c1 */
            {8'h00}, /* 0x06c0 */
            {8'h00}, /* 0x06bf */
            {8'h00}, /* 0x06be */
            {8'h00}, /* 0x06bd */
            {8'h00}, /* 0x06bc */
            {8'h00}, /* 0x06bb */
            {8'h00}, /* 0x06ba */
            {8'h00}, /* 0x06b9 */
            {8'h00}, /* 0x06b8 */
            {8'h00}, /* 0x06b7 */
            {8'h00}, /* 0x06b6 */
            {8'h00}, /* 0x06b5 */
            {8'h00}, /* 0x06b4 */
            {8'h00}, /* 0x06b3 */
            {8'h00}, /* 0x06b2 */
            {8'h00}, /* 0x06b1 */
            {8'h00}, /* 0x06b0 */
            {8'h00}, /* 0x06af */
            {8'h00}, /* 0x06ae */
            {8'h00}, /* 0x06ad */
            {8'h00}, /* 0x06ac */
            {8'h00}, /* 0x06ab */
            {8'h00}, /* 0x06aa */
            {8'h00}, /* 0x06a9 */
            {8'h00}, /* 0x06a8 */
            {8'h00}, /* 0x06a7 */
            {8'h00}, /* 0x06a6 */
            {8'h00}, /* 0x06a5 */
            {8'h00}, /* 0x06a4 */
            {8'h00}, /* 0x06a3 */
            {8'h00}, /* 0x06a2 */
            {8'h00}, /* 0x06a1 */
            {8'h00}, /* 0x06a0 */
            {8'h00}, /* 0x069f */
            {8'h00}, /* 0x069e */
            {8'h00}, /* 0x069d */
            {8'h00}, /* 0x069c */
            {8'h00}, /* 0x069b */
            {8'h00}, /* 0x069a */
            {8'h00}, /* 0x0699 */
            {8'h00}, /* 0x0698 */
            {8'h00}, /* 0x0697 */
            {8'h00}, /* 0x0696 */
            {8'h00}, /* 0x0695 */
            {8'h00}, /* 0x0694 */
            {8'h00}, /* 0x0693 */
            {8'h00}, /* 0x0692 */
            {8'h00}, /* 0x0691 */
            {8'h00}, /* 0x0690 */
            {8'h00}, /* 0x068f */
            {8'h00}, /* 0x068e */
            {8'h00}, /* 0x068d */
            {8'h00}, /* 0x068c */
            {8'h00}, /* 0x068b */
            {8'h00}, /* 0x068a */
            {8'h00}, /* 0x0689 */
            {8'h00}, /* 0x0688 */
            {8'h00}, /* 0x0687 */
            {8'h00}, /* 0x0686 */
            {8'h00}, /* 0x0685 */
            {8'h00}, /* 0x0684 */
            {8'h00}, /* 0x0683 */
            {8'h00}, /* 0x0682 */
            {8'h00}, /* 0x0681 */
            {8'h00}, /* 0x0680 */
            {8'h00}, /* 0x067f */
            {8'h00}, /* 0x067e */
            {8'h00}, /* 0x067d */
            {8'h00}, /* 0x067c */
            {8'h00}, /* 0x067b */
            {8'h00}, /* 0x067a */
            {8'h00}, /* 0x0679 */
            {8'h00}, /* 0x0678 */
            {8'h00}, /* 0x0677 */
            {8'h00}, /* 0x0676 */
            {8'h00}, /* 0x0675 */
            {8'h00}, /* 0x0674 */
            {8'h00}, /* 0x0673 */
            {8'h00}, /* 0x0672 */
            {8'h00}, /* 0x0671 */
            {8'h00}, /* 0x0670 */
            {8'h00}, /* 0x066f */
            {8'h00}, /* 0x066e */
            {8'h00}, /* 0x066d */
            {8'h00}, /* 0x066c */
            {8'h00}, /* 0x066b */
            {8'h00}, /* 0x066a */
            {8'h00}, /* 0x0669 */
            {8'h00}, /* 0x0668 */
            {8'h00}, /* 0x0667 */
            {8'h00}, /* 0x0666 */
            {8'h00}, /* 0x0665 */
            {8'h00}, /* 0x0664 */
            {8'h00}, /* 0x0663 */
            {8'h00}, /* 0x0662 */
            {8'h00}, /* 0x0661 */
            {8'h00}, /* 0x0660 */
            {8'h00}, /* 0x065f */
            {8'h00}, /* 0x065e */
            {8'h00}, /* 0x065d */
            {8'h00}, /* 0x065c */
            {8'h00}, /* 0x065b */
            {8'h00}, /* 0x065a */
            {8'h00}, /* 0x0659 */
            {8'h00}, /* 0x0658 */
            {8'h00}, /* 0x0657 */
            {8'h00}, /* 0x0656 */
            {8'h00}, /* 0x0655 */
            {8'h00}, /* 0x0654 */
            {8'h00}, /* 0x0653 */
            {8'h00}, /* 0x0652 */
            {8'h00}, /* 0x0651 */
            {8'h00}, /* 0x0650 */
            {8'h00}, /* 0x064f */
            {8'h00}, /* 0x064e */
            {8'h00}, /* 0x064d */
            {8'h00}, /* 0x064c */
            {8'h00}, /* 0x064b */
            {8'h00}, /* 0x064a */
            {8'h00}, /* 0x0649 */
            {8'h00}, /* 0x0648 */
            {8'h00}, /* 0x0647 */
            {8'h00}, /* 0x0646 */
            {8'h00}, /* 0x0645 */
            {8'h00}, /* 0x0644 */
            {8'h00}, /* 0x0643 */
            {8'h00}, /* 0x0642 */
            {8'h00}, /* 0x0641 */
            {8'h00}, /* 0x0640 */
            {8'h00}, /* 0x063f */
            {8'h00}, /* 0x063e */
            {8'h00}, /* 0x063d */
            {8'h00}, /* 0x063c */
            {8'h00}, /* 0x063b */
            {8'h00}, /* 0x063a */
            {8'h00}, /* 0x0639 */
            {8'h00}, /* 0x0638 */
            {8'h00}, /* 0x0637 */
            {8'h00}, /* 0x0636 */
            {8'h00}, /* 0x0635 */
            {8'h00}, /* 0x0634 */
            {8'h00}, /* 0x0633 */
            {8'h00}, /* 0x0632 */
            {8'h00}, /* 0x0631 */
            {8'h00}, /* 0x0630 */
            {8'h00}, /* 0x062f */
            {8'h00}, /* 0x062e */
            {8'h00}, /* 0x062d */
            {8'h00}, /* 0x062c */
            {8'h00}, /* 0x062b */
            {8'h00}, /* 0x062a */
            {8'h00}, /* 0x0629 */
            {8'h00}, /* 0x0628 */
            {8'h00}, /* 0x0627 */
            {8'h00}, /* 0x0626 */
            {8'h00}, /* 0x0625 */
            {8'h00}, /* 0x0624 */
            {8'h00}, /* 0x0623 */
            {8'h00}, /* 0x0622 */
            {8'h00}, /* 0x0621 */
            {8'h00}, /* 0x0620 */
            {8'h00}, /* 0x061f */
            {8'h00}, /* 0x061e */
            {8'h00}, /* 0x061d */
            {8'h00}, /* 0x061c */
            {8'h00}, /* 0x061b */
            {8'h00}, /* 0x061a */
            {8'h00}, /* 0x0619 */
            {8'h00}, /* 0x0618 */
            {8'h00}, /* 0x0617 */
            {8'h00}, /* 0x0616 */
            {8'h00}, /* 0x0615 */
            {8'h00}, /* 0x0614 */
            {8'h00}, /* 0x0613 */
            {8'h00}, /* 0x0612 */
            {8'h00}, /* 0x0611 */
            {8'h00}, /* 0x0610 */
            {8'h00}, /* 0x060f */
            {8'h00}, /* 0x060e */
            {8'h00}, /* 0x060d */
            {8'h00}, /* 0x060c */
            {8'h00}, /* 0x060b */
            {8'h00}, /* 0x060a */
            {8'h00}, /* 0x0609 */
            {8'h00}, /* 0x0608 */
            {8'h00}, /* 0x0607 */
            {8'h00}, /* 0x0606 */
            {8'h00}, /* 0x0605 */
            {8'h00}, /* 0x0604 */
            {8'h00}, /* 0x0603 */
            {8'h00}, /* 0x0602 */
            {8'h00}, /* 0x0601 */
            {8'h00}, /* 0x0600 */
            {8'h00}, /* 0x05ff */
            {8'h00}, /* 0x05fe */
            {8'h00}, /* 0x05fd */
            {8'h00}, /* 0x05fc */
            {8'h00}, /* 0x05fb */
            {8'h00}, /* 0x05fa */
            {8'h00}, /* 0x05f9 */
            {8'h00}, /* 0x05f8 */
            {8'h00}, /* 0x05f7 */
            {8'h00}, /* 0x05f6 */
            {8'h00}, /* 0x05f5 */
            {8'h00}, /* 0x05f4 */
            {8'h00}, /* 0x05f3 */
            {8'h00}, /* 0x05f2 */
            {8'h00}, /* 0x05f1 */
            {8'h00}, /* 0x05f0 */
            {8'h00}, /* 0x05ef */
            {8'h00}, /* 0x05ee */
            {8'h00}, /* 0x05ed */
            {8'h00}, /* 0x05ec */
            {8'h00}, /* 0x05eb */
            {8'h00}, /* 0x05ea */
            {8'h00}, /* 0x05e9 */
            {8'h00}, /* 0x05e8 */
            {8'h00}, /* 0x05e7 */
            {8'h00}, /* 0x05e6 */
            {8'h00}, /* 0x05e5 */
            {8'h00}, /* 0x05e4 */
            {8'h00}, /* 0x05e3 */
            {8'h00}, /* 0x05e2 */
            {8'h00}, /* 0x05e1 */
            {8'h00}, /* 0x05e0 */
            {8'h00}, /* 0x05df */
            {8'h00}, /* 0x05de */
            {8'h00}, /* 0x05dd */
            {8'h00}, /* 0x05dc */
            {8'h00}, /* 0x05db */
            {8'h00}, /* 0x05da */
            {8'h00}, /* 0x05d9 */
            {8'h00}, /* 0x05d8 */
            {8'h00}, /* 0x05d7 */
            {8'h00}, /* 0x05d6 */
            {8'h00}, /* 0x05d5 */
            {8'h00}, /* 0x05d4 */
            {8'h00}, /* 0x05d3 */
            {8'h00}, /* 0x05d2 */
            {8'h00}, /* 0x05d1 */
            {8'h00}, /* 0x05d0 */
            {8'h00}, /* 0x05cf */
            {8'h00}, /* 0x05ce */
            {8'h00}, /* 0x05cd */
            {8'h00}, /* 0x05cc */
            {8'h00}, /* 0x05cb */
            {8'h00}, /* 0x05ca */
            {8'h00}, /* 0x05c9 */
            {8'h00}, /* 0x05c8 */
            {8'h00}, /* 0x05c7 */
            {8'h00}, /* 0x05c6 */
            {8'h00}, /* 0x05c5 */
            {8'h00}, /* 0x05c4 */
            {8'h00}, /* 0x05c3 */
            {8'h00}, /* 0x05c2 */
            {8'h00}, /* 0x05c1 */
            {8'h00}, /* 0x05c0 */
            {8'h00}, /* 0x05bf */
            {8'h00}, /* 0x05be */
            {8'h00}, /* 0x05bd */
            {8'h00}, /* 0x05bc */
            {8'h00}, /* 0x05bb */
            {8'h00}, /* 0x05ba */
            {8'h00}, /* 0x05b9 */
            {8'h00}, /* 0x05b8 */
            {8'h00}, /* 0x05b7 */
            {8'h00}, /* 0x05b6 */
            {8'h00}, /* 0x05b5 */
            {8'h00}, /* 0x05b4 */
            {8'h00}, /* 0x05b3 */
            {8'h00}, /* 0x05b2 */
            {8'h00}, /* 0x05b1 */
            {8'h00}, /* 0x05b0 */
            {8'h00}, /* 0x05af */
            {8'h00}, /* 0x05ae */
            {8'h00}, /* 0x05ad */
            {8'h00}, /* 0x05ac */
            {8'h00}, /* 0x05ab */
            {8'h00}, /* 0x05aa */
            {8'h00}, /* 0x05a9 */
            {8'h00}, /* 0x05a8 */
            {8'h00}, /* 0x05a7 */
            {8'h00}, /* 0x05a6 */
            {8'h00}, /* 0x05a5 */
            {8'h00}, /* 0x05a4 */
            {8'h00}, /* 0x05a3 */
            {8'h00}, /* 0x05a2 */
            {8'h00}, /* 0x05a1 */
            {8'h00}, /* 0x05a0 */
            {8'h00}, /* 0x059f */
            {8'h00}, /* 0x059e */
            {8'h00}, /* 0x059d */
            {8'h00}, /* 0x059c */
            {8'h00}, /* 0x059b */
            {8'h00}, /* 0x059a */
            {8'h00}, /* 0x0599 */
            {8'h00}, /* 0x0598 */
            {8'h00}, /* 0x0597 */
            {8'h00}, /* 0x0596 */
            {8'h00}, /* 0x0595 */
            {8'h00}, /* 0x0594 */
            {8'h00}, /* 0x0593 */
            {8'h00}, /* 0x0592 */
            {8'h00}, /* 0x0591 */
            {8'h00}, /* 0x0590 */
            {8'h00}, /* 0x058f */
            {8'h00}, /* 0x058e */
            {8'h00}, /* 0x058d */
            {8'h00}, /* 0x058c */
            {8'h00}, /* 0x058b */
            {8'h00}, /* 0x058a */
            {8'h00}, /* 0x0589 */
            {8'h00}, /* 0x0588 */
            {8'h00}, /* 0x0587 */
            {8'h00}, /* 0x0586 */
            {8'h00}, /* 0x0585 */
            {8'h00}, /* 0x0584 */
            {8'h00}, /* 0x0583 */
            {8'h00}, /* 0x0582 */
            {8'h00}, /* 0x0581 */
            {8'h00}, /* 0x0580 */
            {8'h00}, /* 0x057f */
            {8'h00}, /* 0x057e */
            {8'h00}, /* 0x057d */
            {8'h00}, /* 0x057c */
            {8'h00}, /* 0x057b */
            {8'h00}, /* 0x057a */
            {8'h00}, /* 0x0579 */
            {8'h00}, /* 0x0578 */
            {8'h00}, /* 0x0577 */
            {8'h00}, /* 0x0576 */
            {8'h00}, /* 0x0575 */
            {8'h00}, /* 0x0574 */
            {8'h00}, /* 0x0573 */
            {8'h00}, /* 0x0572 */
            {8'h00}, /* 0x0571 */
            {8'h00}, /* 0x0570 */
            {8'h00}, /* 0x056f */
            {8'h00}, /* 0x056e */
            {8'h00}, /* 0x056d */
            {8'h00}, /* 0x056c */
            {8'h00}, /* 0x056b */
            {8'h00}, /* 0x056a */
            {8'h00}, /* 0x0569 */
            {8'h00}, /* 0x0568 */
            {8'h00}, /* 0x0567 */
            {8'h00}, /* 0x0566 */
            {8'h00}, /* 0x0565 */
            {8'h00}, /* 0x0564 */
            {8'h00}, /* 0x0563 */
            {8'h00}, /* 0x0562 */
            {8'h00}, /* 0x0561 */
            {8'h00}, /* 0x0560 */
            {8'h00}, /* 0x055f */
            {8'h00}, /* 0x055e */
            {8'h00}, /* 0x055d */
            {8'h00}, /* 0x055c */
            {8'h00}, /* 0x055b */
            {8'h00}, /* 0x055a */
            {8'h00}, /* 0x0559 */
            {8'h00}, /* 0x0558 */
            {8'h00}, /* 0x0557 */
            {8'h00}, /* 0x0556 */
            {8'h00}, /* 0x0555 */
            {8'h00}, /* 0x0554 */
            {8'h00}, /* 0x0553 */
            {8'h00}, /* 0x0552 */
            {8'h00}, /* 0x0551 */
            {8'h00}, /* 0x0550 */
            {8'h00}, /* 0x054f */
            {8'h00}, /* 0x054e */
            {8'h00}, /* 0x054d */
            {8'h00}, /* 0x054c */
            {8'h00}, /* 0x054b */
            {8'h00}, /* 0x054a */
            {8'h00}, /* 0x0549 */
            {8'h00}, /* 0x0548 */
            {8'h00}, /* 0x0547 */
            {8'h00}, /* 0x0546 */
            {8'h00}, /* 0x0545 */
            {8'h00}, /* 0x0544 */
            {8'h00}, /* 0x0543 */
            {8'h00}, /* 0x0542 */
            {8'h00}, /* 0x0541 */
            {8'h00}, /* 0x0540 */
            {8'h00}, /* 0x053f */
            {8'h00}, /* 0x053e */
            {8'h00}, /* 0x053d */
            {8'h00}, /* 0x053c */
            {8'h00}, /* 0x053b */
            {8'h00}, /* 0x053a */
            {8'h00}, /* 0x0539 */
            {8'h00}, /* 0x0538 */
            {8'h00}, /* 0x0537 */
            {8'h00}, /* 0x0536 */
            {8'h00}, /* 0x0535 */
            {8'h00}, /* 0x0534 */
            {8'h00}, /* 0x0533 */
            {8'h00}, /* 0x0532 */
            {8'h00}, /* 0x0531 */
            {8'h00}, /* 0x0530 */
            {8'h00}, /* 0x052f */
            {8'h00}, /* 0x052e */
            {8'h00}, /* 0x052d */
            {8'h00}, /* 0x052c */
            {8'h00}, /* 0x052b */
            {8'h00}, /* 0x052a */
            {8'h00}, /* 0x0529 */
            {8'h00}, /* 0x0528 */
            {8'h00}, /* 0x0527 */
            {8'h00}, /* 0x0526 */
            {8'h00}, /* 0x0525 */
            {8'h00}, /* 0x0524 */
            {8'h00}, /* 0x0523 */
            {8'h00}, /* 0x0522 */
            {8'h00}, /* 0x0521 */
            {8'h00}, /* 0x0520 */
            {8'h00}, /* 0x051f */
            {8'h00}, /* 0x051e */
            {8'h00}, /* 0x051d */
            {8'h00}, /* 0x051c */
            {8'h00}, /* 0x051b */
            {8'h00}, /* 0x051a */
            {8'h00}, /* 0x0519 */
            {8'h00}, /* 0x0518 */
            {8'h00}, /* 0x0517 */
            {8'h00}, /* 0x0516 */
            {8'h00}, /* 0x0515 */
            {8'h00}, /* 0x0514 */
            {8'h00}, /* 0x0513 */
            {8'h00}, /* 0x0512 */
            {8'h00}, /* 0x0511 */
            {8'h00}, /* 0x0510 */
            {8'h00}, /* 0x050f */
            {8'h00}, /* 0x050e */
            {8'h00}, /* 0x050d */
            {8'h00}, /* 0x050c */
            {8'h00}, /* 0x050b */
            {8'h00}, /* 0x050a */
            {8'h00}, /* 0x0509 */
            {8'h00}, /* 0x0508 */
            {8'h00}, /* 0x0507 */
            {8'h00}, /* 0x0506 */
            {8'h00}, /* 0x0505 */
            {8'h00}, /* 0x0504 */
            {8'h00}, /* 0x0503 */
            {8'h00}, /* 0x0502 */
            {8'h00}, /* 0x0501 */
            {8'h00}, /* 0x0500 */
            {8'h00}, /* 0x04ff */
            {8'h00}, /* 0x04fe */
            {8'h00}, /* 0x04fd */
            {8'h00}, /* 0x04fc */
            {8'h00}, /* 0x04fb */
            {8'h00}, /* 0x04fa */
            {8'h00}, /* 0x04f9 */
            {8'h00}, /* 0x04f8 */
            {8'h00}, /* 0x04f7 */
            {8'h00}, /* 0x04f6 */
            {8'h00}, /* 0x04f5 */
            {8'h00}, /* 0x04f4 */
            {8'h00}, /* 0x04f3 */
            {8'h00}, /* 0x04f2 */
            {8'h00}, /* 0x04f1 */
            {8'h00}, /* 0x04f0 */
            {8'h00}, /* 0x04ef */
            {8'h00}, /* 0x04ee */
            {8'h00}, /* 0x04ed */
            {8'h00}, /* 0x04ec */
            {8'h00}, /* 0x04eb */
            {8'h00}, /* 0x04ea */
            {8'h00}, /* 0x04e9 */
            {8'h00}, /* 0x04e8 */
            {8'h00}, /* 0x04e7 */
            {8'h00}, /* 0x04e6 */
            {8'h00}, /* 0x04e5 */
            {8'h00}, /* 0x04e4 */
            {8'h00}, /* 0x04e3 */
            {8'h00}, /* 0x04e2 */
            {8'h00}, /* 0x04e1 */
            {8'h00}, /* 0x04e0 */
            {8'h00}, /* 0x04df */
            {8'h00}, /* 0x04de */
            {8'h00}, /* 0x04dd */
            {8'h00}, /* 0x04dc */
            {8'h00}, /* 0x04db */
            {8'h00}, /* 0x04da */
            {8'h00}, /* 0x04d9 */
            {8'h00}, /* 0x04d8 */
            {8'h00}, /* 0x04d7 */
            {8'h00}, /* 0x04d6 */
            {8'h00}, /* 0x04d5 */
            {8'h00}, /* 0x04d4 */
            {8'h00}, /* 0x04d3 */
            {8'h00}, /* 0x04d2 */
            {8'h00}, /* 0x04d1 */
            {8'h00}, /* 0x04d0 */
            {8'h00}, /* 0x04cf */
            {8'h00}, /* 0x04ce */
            {8'h00}, /* 0x04cd */
            {8'h00}, /* 0x04cc */
            {8'h00}, /* 0x04cb */
            {8'h00}, /* 0x04ca */
            {8'h00}, /* 0x04c9 */
            {8'h00}, /* 0x04c8 */
            {8'h00}, /* 0x04c7 */
            {8'h00}, /* 0x04c6 */
            {8'h00}, /* 0x04c5 */
            {8'h00}, /* 0x04c4 */
            {8'h00}, /* 0x04c3 */
            {8'h00}, /* 0x04c2 */
            {8'h00}, /* 0x04c1 */
            {8'h00}, /* 0x04c0 */
            {8'h00}, /* 0x04bf */
            {8'h00}, /* 0x04be */
            {8'h00}, /* 0x04bd */
            {8'h00}, /* 0x04bc */
            {8'h00}, /* 0x04bb */
            {8'h00}, /* 0x04ba */
            {8'h00}, /* 0x04b9 */
            {8'h00}, /* 0x04b8 */
            {8'h00}, /* 0x04b7 */
            {8'h00}, /* 0x04b6 */
            {8'h00}, /* 0x04b5 */
            {8'h00}, /* 0x04b4 */
            {8'h00}, /* 0x04b3 */
            {8'h00}, /* 0x04b2 */
            {8'h00}, /* 0x04b1 */
            {8'h00}, /* 0x04b0 */
            {8'h00}, /* 0x04af */
            {8'h00}, /* 0x04ae */
            {8'h00}, /* 0x04ad */
            {8'h00}, /* 0x04ac */
            {8'h00}, /* 0x04ab */
            {8'h00}, /* 0x04aa */
            {8'h00}, /* 0x04a9 */
            {8'h00}, /* 0x04a8 */
            {8'h00}, /* 0x04a7 */
            {8'h00}, /* 0x04a6 */
            {8'h00}, /* 0x04a5 */
            {8'h00}, /* 0x04a4 */
            {8'h00}, /* 0x04a3 */
            {8'h00}, /* 0x04a2 */
            {8'h00}, /* 0x04a1 */
            {8'h00}, /* 0x04a0 */
            {8'h00}, /* 0x049f */
            {8'h00}, /* 0x049e */
            {8'h00}, /* 0x049d */
            {8'h00}, /* 0x049c */
            {8'h00}, /* 0x049b */
            {8'h00}, /* 0x049a */
            {8'h00}, /* 0x0499 */
            {8'h00}, /* 0x0498 */
            {8'h00}, /* 0x0497 */
            {8'h00}, /* 0x0496 */
            {8'h00}, /* 0x0495 */
            {8'h00}, /* 0x0494 */
            {8'h00}, /* 0x0493 */
            {8'h00}, /* 0x0492 */
            {8'h00}, /* 0x0491 */
            {8'h00}, /* 0x0490 */
            {8'h00}, /* 0x048f */
            {8'h00}, /* 0x048e */
            {8'h00}, /* 0x048d */
            {8'h00}, /* 0x048c */
            {8'h00}, /* 0x048b */
            {8'h00}, /* 0x048a */
            {8'h00}, /* 0x0489 */
            {8'h00}, /* 0x0488 */
            {8'h00}, /* 0x0487 */
            {8'h00}, /* 0x0486 */
            {8'h00}, /* 0x0485 */
            {8'h00}, /* 0x0484 */
            {8'h00}, /* 0x0483 */
            {8'h00}, /* 0x0482 */
            {8'h00}, /* 0x0481 */
            {8'h00}, /* 0x0480 */
            {8'h00}, /* 0x047f */
            {8'h00}, /* 0x047e */
            {8'h00}, /* 0x047d */
            {8'h00}, /* 0x047c */
            {8'h00}, /* 0x047b */
            {8'h00}, /* 0x047a */
            {8'h00}, /* 0x0479 */
            {8'h00}, /* 0x0478 */
            {8'h00}, /* 0x0477 */
            {8'h00}, /* 0x0476 */
            {8'h00}, /* 0x0475 */
            {8'h00}, /* 0x0474 */
            {8'h00}, /* 0x0473 */
            {8'h00}, /* 0x0472 */
            {8'h00}, /* 0x0471 */
            {8'h00}, /* 0x0470 */
            {8'h00}, /* 0x046f */
            {8'h00}, /* 0x046e */
            {8'h00}, /* 0x046d */
            {8'h00}, /* 0x046c */
            {8'h00}, /* 0x046b */
            {8'h00}, /* 0x046a */
            {8'h00}, /* 0x0469 */
            {8'h00}, /* 0x0468 */
            {8'h00}, /* 0x0467 */
            {8'h00}, /* 0x0466 */
            {8'h00}, /* 0x0465 */
            {8'h00}, /* 0x0464 */
            {8'h00}, /* 0x0463 */
            {8'h00}, /* 0x0462 */
            {8'h00}, /* 0x0461 */
            {8'h00}, /* 0x0460 */
            {8'h00}, /* 0x045f */
            {8'h00}, /* 0x045e */
            {8'h00}, /* 0x045d */
            {8'h00}, /* 0x045c */
            {8'h00}, /* 0x045b */
            {8'h00}, /* 0x045a */
            {8'h00}, /* 0x0459 */
            {8'h00}, /* 0x0458 */
            {8'h00}, /* 0x0457 */
            {8'h00}, /* 0x0456 */
            {8'h00}, /* 0x0455 */
            {8'h00}, /* 0x0454 */
            {8'h00}, /* 0x0453 */
            {8'h00}, /* 0x0452 */
            {8'h00}, /* 0x0451 */
            {8'h00}, /* 0x0450 */
            {8'h00}, /* 0x044f */
            {8'h00}, /* 0x044e */
            {8'h00}, /* 0x044d */
            {8'h00}, /* 0x044c */
            {8'h00}, /* 0x044b */
            {8'h00}, /* 0x044a */
            {8'h00}, /* 0x0449 */
            {8'h00}, /* 0x0448 */
            {8'h00}, /* 0x0447 */
            {8'h00}, /* 0x0446 */
            {8'h00}, /* 0x0445 */
            {8'h00}, /* 0x0444 */
            {8'h00}, /* 0x0443 */
            {8'h00}, /* 0x0442 */
            {8'h00}, /* 0x0441 */
            {8'h00}, /* 0x0440 */
            {8'h00}, /* 0x043f */
            {8'h00}, /* 0x043e */
            {8'h00}, /* 0x043d */
            {8'h00}, /* 0x043c */
            {8'h00}, /* 0x043b */
            {8'h00}, /* 0x043a */
            {8'h00}, /* 0x0439 */
            {8'h00}, /* 0x0438 */
            {8'h00}, /* 0x0437 */
            {8'h00}, /* 0x0436 */
            {8'h00}, /* 0x0435 */
            {8'h00}, /* 0x0434 */
            {8'h00}, /* 0x0433 */
            {8'h00}, /* 0x0432 */
            {8'h00}, /* 0x0431 */
            {8'h00}, /* 0x0430 */
            {8'h00}, /* 0x042f */
            {8'h00}, /* 0x042e */
            {8'h00}, /* 0x042d */
            {8'h00}, /* 0x042c */
            {8'h00}, /* 0x042b */
            {8'h00}, /* 0x042a */
            {8'h00}, /* 0x0429 */
            {8'h00}, /* 0x0428 */
            {8'h00}, /* 0x0427 */
            {8'h00}, /* 0x0426 */
            {8'h00}, /* 0x0425 */
            {8'h00}, /* 0x0424 */
            {8'h00}, /* 0x0423 */
            {8'h00}, /* 0x0422 */
            {8'h00}, /* 0x0421 */
            {8'h00}, /* 0x0420 */
            {8'h00}, /* 0x041f */
            {8'h00}, /* 0x041e */
            {8'h00}, /* 0x041d */
            {8'h00}, /* 0x041c */
            {8'h00}, /* 0x041b */
            {8'h00}, /* 0x041a */
            {8'h00}, /* 0x0419 */
            {8'h00}, /* 0x0418 */
            {8'h00}, /* 0x0417 */
            {8'h00}, /* 0x0416 */
            {8'h00}, /* 0x0415 */
            {8'h00}, /* 0x0414 */
            {8'h00}, /* 0x0413 */
            {8'h00}, /* 0x0412 */
            {8'h00}, /* 0x0411 */
            {8'h00}, /* 0x0410 */
            {8'h00}, /* 0x040f */
            {8'h00}, /* 0x040e */
            {8'h00}, /* 0x040d */
            {8'h00}, /* 0x040c */
            {8'h00}, /* 0x040b */
            {8'h00}, /* 0x040a */
            {8'h00}, /* 0x0409 */
            {8'h00}, /* 0x0408 */
            {8'h00}, /* 0x0407 */
            {8'h00}, /* 0x0406 */
            {8'h00}, /* 0x0405 */
            {8'h00}, /* 0x0404 */
            {8'h00}, /* 0x0403 */
            {8'h00}, /* 0x0402 */
            {8'h00}, /* 0x0401 */
            {8'h00}, /* 0x0400 */
            {8'h00}, /* 0x03ff */
            {8'h00}, /* 0x03fe */
            {8'h00}, /* 0x03fd */
            {8'h00}, /* 0x03fc */
            {8'h00}, /* 0x03fb */
            {8'h00}, /* 0x03fa */
            {8'h00}, /* 0x03f9 */
            {8'h00}, /* 0x03f8 */
            {8'h00}, /* 0x03f7 */
            {8'h00}, /* 0x03f6 */
            {8'h00}, /* 0x03f5 */
            {8'h00}, /* 0x03f4 */
            {8'h00}, /* 0x03f3 */
            {8'h00}, /* 0x03f2 */
            {8'h00}, /* 0x03f1 */
            {8'h00}, /* 0x03f0 */
            {8'h00}, /* 0x03ef */
            {8'h00}, /* 0x03ee */
            {8'h00}, /* 0x03ed */
            {8'h00}, /* 0x03ec */
            {8'h00}, /* 0x03eb */
            {8'h00}, /* 0x03ea */
            {8'h00}, /* 0x03e9 */
            {8'h00}, /* 0x03e8 */
            {8'h00}, /* 0x03e7 */
            {8'h00}, /* 0x03e6 */
            {8'h00}, /* 0x03e5 */
            {8'h00}, /* 0x03e4 */
            {8'h00}, /* 0x03e3 */
            {8'h00}, /* 0x03e2 */
            {8'h00}, /* 0x03e1 */
            {8'h00}, /* 0x03e0 */
            {8'h00}, /* 0x03df */
            {8'h00}, /* 0x03de */
            {8'h00}, /* 0x03dd */
            {8'h00}, /* 0x03dc */
            {8'h00}, /* 0x03db */
            {8'h00}, /* 0x03da */
            {8'h00}, /* 0x03d9 */
            {8'h00}, /* 0x03d8 */
            {8'h00}, /* 0x03d7 */
            {8'h00}, /* 0x03d6 */
            {8'h00}, /* 0x03d5 */
            {8'h00}, /* 0x03d4 */
            {8'h00}, /* 0x03d3 */
            {8'h00}, /* 0x03d2 */
            {8'h00}, /* 0x03d1 */
            {8'h00}, /* 0x03d0 */
            {8'h00}, /* 0x03cf */
            {8'h00}, /* 0x03ce */
            {8'h00}, /* 0x03cd */
            {8'h00}, /* 0x03cc */
            {8'h00}, /* 0x03cb */
            {8'h00}, /* 0x03ca */
            {8'h00}, /* 0x03c9 */
            {8'h00}, /* 0x03c8 */
            {8'h00}, /* 0x03c7 */
            {8'h00}, /* 0x03c6 */
            {8'h00}, /* 0x03c5 */
            {8'h00}, /* 0x03c4 */
            {8'h00}, /* 0x03c3 */
            {8'h00}, /* 0x03c2 */
            {8'h00}, /* 0x03c1 */
            {8'h00}, /* 0x03c0 */
            {8'h00}, /* 0x03bf */
            {8'h00}, /* 0x03be */
            {8'h00}, /* 0x03bd */
            {8'h00}, /* 0x03bc */
            {8'h00}, /* 0x03bb */
            {8'h00}, /* 0x03ba */
            {8'h00}, /* 0x03b9 */
            {8'h00}, /* 0x03b8 */
            {8'h00}, /* 0x03b7 */
            {8'h00}, /* 0x03b6 */
            {8'h00}, /* 0x03b5 */
            {8'h00}, /* 0x03b4 */
            {8'h00}, /* 0x03b3 */
            {8'h00}, /* 0x03b2 */
            {8'h00}, /* 0x03b1 */
            {8'h00}, /* 0x03b0 */
            {8'h00}, /* 0x03af */
            {8'h00}, /* 0x03ae */
            {8'h00}, /* 0x03ad */
            {8'h00}, /* 0x03ac */
            {8'h00}, /* 0x03ab */
            {8'h00}, /* 0x03aa */
            {8'h00}, /* 0x03a9 */
            {8'h00}, /* 0x03a8 */
            {8'h00}, /* 0x03a7 */
            {8'h00}, /* 0x03a6 */
            {8'h00}, /* 0x03a5 */
            {8'h00}, /* 0x03a4 */
            {8'h00}, /* 0x03a3 */
            {8'h00}, /* 0x03a2 */
            {8'h00}, /* 0x03a1 */
            {8'h00}, /* 0x03a0 */
            {8'h00}, /* 0x039f */
            {8'h00}, /* 0x039e */
            {8'h00}, /* 0x039d */
            {8'h00}, /* 0x039c */
            {8'h00}, /* 0x039b */
            {8'h00}, /* 0x039a */
            {8'h00}, /* 0x0399 */
            {8'h00}, /* 0x0398 */
            {8'h00}, /* 0x0397 */
            {8'h00}, /* 0x0396 */
            {8'h00}, /* 0x0395 */
            {8'h00}, /* 0x0394 */
            {8'h00}, /* 0x0393 */
            {8'h00}, /* 0x0392 */
            {8'h00}, /* 0x0391 */
            {8'h00}, /* 0x0390 */
            {8'h00}, /* 0x038f */
            {8'h00}, /* 0x038e */
            {8'h00}, /* 0x038d */
            {8'h00}, /* 0x038c */
            {8'h00}, /* 0x038b */
            {8'h00}, /* 0x038a */
            {8'h00}, /* 0x0389 */
            {8'h00}, /* 0x0388 */
            {8'h00}, /* 0x0387 */
            {8'h00}, /* 0x0386 */
            {8'h00}, /* 0x0385 */
            {8'h00}, /* 0x0384 */
            {8'h00}, /* 0x0383 */
            {8'h00}, /* 0x0382 */
            {8'h00}, /* 0x0381 */
            {8'h00}, /* 0x0380 */
            {8'h00}, /* 0x037f */
            {8'h00}, /* 0x037e */
            {8'h00}, /* 0x037d */
            {8'h00}, /* 0x037c */
            {8'h00}, /* 0x037b */
            {8'h00}, /* 0x037a */
            {8'h00}, /* 0x0379 */
            {8'h00}, /* 0x0378 */
            {8'h00}, /* 0x0377 */
            {8'h00}, /* 0x0376 */
            {8'h00}, /* 0x0375 */
            {8'h00}, /* 0x0374 */
            {8'h00}, /* 0x0373 */
            {8'h00}, /* 0x0372 */
            {8'h00}, /* 0x0371 */
            {8'h00}, /* 0x0370 */
            {8'h00}, /* 0x036f */
            {8'h00}, /* 0x036e */
            {8'h00}, /* 0x036d */
            {8'h00}, /* 0x036c */
            {8'h00}, /* 0x036b */
            {8'h00}, /* 0x036a */
            {8'h00}, /* 0x0369 */
            {8'h00}, /* 0x0368 */
            {8'h00}, /* 0x0367 */
            {8'h00}, /* 0x0366 */
            {8'h00}, /* 0x0365 */
            {8'h00}, /* 0x0364 */
            {8'h00}, /* 0x0363 */
            {8'h00}, /* 0x0362 */
            {8'h00}, /* 0x0361 */
            {8'h00}, /* 0x0360 */
            {8'h00}, /* 0x035f */
            {8'h00}, /* 0x035e */
            {8'h00}, /* 0x035d */
            {8'h00}, /* 0x035c */
            {8'h00}, /* 0x035b */
            {8'h00}, /* 0x035a */
            {8'h00}, /* 0x0359 */
            {8'h00}, /* 0x0358 */
            {8'h00}, /* 0x0357 */
            {8'h00}, /* 0x0356 */
            {8'h00}, /* 0x0355 */
            {8'h00}, /* 0x0354 */
            {8'h00}, /* 0x0353 */
            {8'h00}, /* 0x0352 */
            {8'h00}, /* 0x0351 */
            {8'h00}, /* 0x0350 */
            {8'h00}, /* 0x034f */
            {8'h00}, /* 0x034e */
            {8'h00}, /* 0x034d */
            {8'h00}, /* 0x034c */
            {8'h00}, /* 0x034b */
            {8'h00}, /* 0x034a */
            {8'h00}, /* 0x0349 */
            {8'h00}, /* 0x0348 */
            {8'h00}, /* 0x0347 */
            {8'h00}, /* 0x0346 */
            {8'h00}, /* 0x0345 */
            {8'h00}, /* 0x0344 */
            {8'h00}, /* 0x0343 */
            {8'h00}, /* 0x0342 */
            {8'h00}, /* 0x0341 */
            {8'h00}, /* 0x0340 */
            {8'h00}, /* 0x033f */
            {8'h00}, /* 0x033e */
            {8'h00}, /* 0x033d */
            {8'h00}, /* 0x033c */
            {8'h00}, /* 0x033b */
            {8'h00}, /* 0x033a */
            {8'h00}, /* 0x0339 */
            {8'h00}, /* 0x0338 */
            {8'h00}, /* 0x0337 */
            {8'h00}, /* 0x0336 */
            {8'h00}, /* 0x0335 */
            {8'h00}, /* 0x0334 */
            {8'h00}, /* 0x0333 */
            {8'h00}, /* 0x0332 */
            {8'h00}, /* 0x0331 */
            {8'h00}, /* 0x0330 */
            {8'h00}, /* 0x032f */
            {8'h00}, /* 0x032e */
            {8'h00}, /* 0x032d */
            {8'h00}, /* 0x032c */
            {8'h00}, /* 0x032b */
            {8'h00}, /* 0x032a */
            {8'h00}, /* 0x0329 */
            {8'h00}, /* 0x0328 */
            {8'h00}, /* 0x0327 */
            {8'h00}, /* 0x0326 */
            {8'h00}, /* 0x0325 */
            {8'h00}, /* 0x0324 */
            {8'h00}, /* 0x0323 */
            {8'h00}, /* 0x0322 */
            {8'h00}, /* 0x0321 */
            {8'h00}, /* 0x0320 */
            {8'h00}, /* 0x031f */
            {8'h00}, /* 0x031e */
            {8'h00}, /* 0x031d */
            {8'h00}, /* 0x031c */
            {8'h00}, /* 0x031b */
            {8'h00}, /* 0x031a */
            {8'h00}, /* 0x0319 */
            {8'h00}, /* 0x0318 */
            {8'h00}, /* 0x0317 */
            {8'h00}, /* 0x0316 */
            {8'h00}, /* 0x0315 */
            {8'h00}, /* 0x0314 */
            {8'h00}, /* 0x0313 */
            {8'h00}, /* 0x0312 */
            {8'h00}, /* 0x0311 */
            {8'h00}, /* 0x0310 */
            {8'h00}, /* 0x030f */
            {8'h00}, /* 0x030e */
            {8'h00}, /* 0x030d */
            {8'h00}, /* 0x030c */
            {8'h00}, /* 0x030b */
            {8'h00}, /* 0x030a */
            {8'h00}, /* 0x0309 */
            {8'h00}, /* 0x0308 */
            {8'h00}, /* 0x0307 */
            {8'h00}, /* 0x0306 */
            {8'h00}, /* 0x0305 */
            {8'h00}, /* 0x0304 */
            {8'h00}, /* 0x0303 */
            {8'h00}, /* 0x0302 */
            {8'h00}, /* 0x0301 */
            {8'h00}, /* 0x0300 */
            {8'h00}, /* 0x02ff */
            {8'h00}, /* 0x02fe */
            {8'h00}, /* 0x02fd */
            {8'h00}, /* 0x02fc */
            {8'h00}, /* 0x02fb */
            {8'h00}, /* 0x02fa */
            {8'h00}, /* 0x02f9 */
            {8'h00}, /* 0x02f8 */
            {8'h00}, /* 0x02f7 */
            {8'h00}, /* 0x02f6 */
            {8'h00}, /* 0x02f5 */
            {8'h00}, /* 0x02f4 */
            {8'h00}, /* 0x02f3 */
            {8'h00}, /* 0x02f2 */
            {8'h00}, /* 0x02f1 */
            {8'h00}, /* 0x02f0 */
            {8'h00}, /* 0x02ef */
            {8'h00}, /* 0x02ee */
            {8'h00}, /* 0x02ed */
            {8'h00}, /* 0x02ec */
            {8'h00}, /* 0x02eb */
            {8'h00}, /* 0x02ea */
            {8'h00}, /* 0x02e9 */
            {8'h00}, /* 0x02e8 */
            {8'h00}, /* 0x02e7 */
            {8'h00}, /* 0x02e6 */
            {8'h00}, /* 0x02e5 */
            {8'h00}, /* 0x02e4 */
            {8'h00}, /* 0x02e3 */
            {8'h00}, /* 0x02e2 */
            {8'h00}, /* 0x02e1 */
            {8'h00}, /* 0x02e0 */
            {8'h00}, /* 0x02df */
            {8'h00}, /* 0x02de */
            {8'h00}, /* 0x02dd */
            {8'h00}, /* 0x02dc */
            {8'h00}, /* 0x02db */
            {8'h00}, /* 0x02da */
            {8'h00}, /* 0x02d9 */
            {8'h00}, /* 0x02d8 */
            {8'h00}, /* 0x02d7 */
            {8'h00}, /* 0x02d6 */
            {8'h00}, /* 0x02d5 */
            {8'h00}, /* 0x02d4 */
            {8'h00}, /* 0x02d3 */
            {8'h00}, /* 0x02d2 */
            {8'h00}, /* 0x02d1 */
            {8'h00}, /* 0x02d0 */
            {8'h00}, /* 0x02cf */
            {8'h00}, /* 0x02ce */
            {8'h00}, /* 0x02cd */
            {8'h00}, /* 0x02cc */
            {8'h00}, /* 0x02cb */
            {8'h00}, /* 0x02ca */
            {8'h00}, /* 0x02c9 */
            {8'h00}, /* 0x02c8 */
            {8'h00}, /* 0x02c7 */
            {8'h00}, /* 0x02c6 */
            {8'h00}, /* 0x02c5 */
            {8'h00}, /* 0x02c4 */
            {8'h00}, /* 0x02c3 */
            {8'h00}, /* 0x02c2 */
            {8'h00}, /* 0x02c1 */
            {8'h00}, /* 0x02c0 */
            {8'h00}, /* 0x02bf */
            {8'h00}, /* 0x02be */
            {8'h00}, /* 0x02bd */
            {8'h00}, /* 0x02bc */
            {8'h00}, /* 0x02bb */
            {8'h00}, /* 0x02ba */
            {8'h00}, /* 0x02b9 */
            {8'h00}, /* 0x02b8 */
            {8'h00}, /* 0x02b7 */
            {8'h00}, /* 0x02b6 */
            {8'h00}, /* 0x02b5 */
            {8'h00}, /* 0x02b4 */
            {8'h00}, /* 0x02b3 */
            {8'h00}, /* 0x02b2 */
            {8'h00}, /* 0x02b1 */
            {8'h00}, /* 0x02b0 */
            {8'h00}, /* 0x02af */
            {8'h00}, /* 0x02ae */
            {8'h00}, /* 0x02ad */
            {8'h00}, /* 0x02ac */
            {8'h00}, /* 0x02ab */
            {8'h00}, /* 0x02aa */
            {8'h00}, /* 0x02a9 */
            {8'h00}, /* 0x02a8 */
            {8'h00}, /* 0x02a7 */
            {8'h00}, /* 0x02a6 */
            {8'h00}, /* 0x02a5 */
            {8'h00}, /* 0x02a4 */
            {8'h00}, /* 0x02a3 */
            {8'h00}, /* 0x02a2 */
            {8'h00}, /* 0x02a1 */
            {8'h00}, /* 0x02a0 */
            {8'h00}, /* 0x029f */
            {8'h00}, /* 0x029e */
            {8'h00}, /* 0x029d */
            {8'h00}, /* 0x029c */
            {8'h00}, /* 0x029b */
            {8'h00}, /* 0x029a */
            {8'h00}, /* 0x0299 */
            {8'h00}, /* 0x0298 */
            {8'h00}, /* 0x0297 */
            {8'h00}, /* 0x0296 */
            {8'h00}, /* 0x0295 */
            {8'h00}, /* 0x0294 */
            {8'h00}, /* 0x0293 */
            {8'h00}, /* 0x0292 */
            {8'h00}, /* 0x0291 */
            {8'h00}, /* 0x0290 */
            {8'h00}, /* 0x028f */
            {8'h00}, /* 0x028e */
            {8'h00}, /* 0x028d */
            {8'h00}, /* 0x028c */
            {8'h00}, /* 0x028b */
            {8'h00}, /* 0x028a */
            {8'h00}, /* 0x0289 */
            {8'h00}, /* 0x0288 */
            {8'h00}, /* 0x0287 */
            {8'h00}, /* 0x0286 */
            {8'h00}, /* 0x0285 */
            {8'h00}, /* 0x0284 */
            {8'h00}, /* 0x0283 */
            {8'h00}, /* 0x0282 */
            {8'h00}, /* 0x0281 */
            {8'h00}, /* 0x0280 */
            {8'h00}, /* 0x027f */
            {8'h00}, /* 0x027e */
            {8'h00}, /* 0x027d */
            {8'h00}, /* 0x027c */
            {8'h00}, /* 0x027b */
            {8'h00}, /* 0x027a */
            {8'h00}, /* 0x0279 */
            {8'h00}, /* 0x0278 */
            {8'h00}, /* 0x0277 */
            {8'h00}, /* 0x0276 */
            {8'h00}, /* 0x0275 */
            {8'h00}, /* 0x0274 */
            {8'h00}, /* 0x0273 */
            {8'h00}, /* 0x0272 */
            {8'h00}, /* 0x0271 */
            {8'h00}, /* 0x0270 */
            {8'h00}, /* 0x026f */
            {8'h00}, /* 0x026e */
            {8'h00}, /* 0x026d */
            {8'h00}, /* 0x026c */
            {8'h00}, /* 0x026b */
            {8'h00}, /* 0x026a */
            {8'h00}, /* 0x0269 */
            {8'h00}, /* 0x0268 */
            {8'h00}, /* 0x0267 */
            {8'h00}, /* 0x0266 */
            {8'h00}, /* 0x0265 */
            {8'h00}, /* 0x0264 */
            {8'h00}, /* 0x0263 */
            {8'h00}, /* 0x0262 */
            {8'h00}, /* 0x0261 */
            {8'h00}, /* 0x0260 */
            {8'h00}, /* 0x025f */
            {8'h00}, /* 0x025e */
            {8'h00}, /* 0x025d */
            {8'h00}, /* 0x025c */
            {8'h00}, /* 0x025b */
            {8'h00}, /* 0x025a */
            {8'h00}, /* 0x0259 */
            {8'h00}, /* 0x0258 */
            {8'h00}, /* 0x0257 */
            {8'h00}, /* 0x0256 */
            {8'h00}, /* 0x0255 */
            {8'h00}, /* 0x0254 */
            {8'h00}, /* 0x0253 */
            {8'h00}, /* 0x0252 */
            {8'h00}, /* 0x0251 */
            {8'h00}, /* 0x0250 */
            {8'h00}, /* 0x024f */
            {8'h00}, /* 0x024e */
            {8'h00}, /* 0x024d */
            {8'h00}, /* 0x024c */
            {8'h00}, /* 0x024b */
            {8'h00}, /* 0x024a */
            {8'h00}, /* 0x0249 */
            {8'h00}, /* 0x0248 */
            {8'h00}, /* 0x0247 */
            {8'h00}, /* 0x0246 */
            {8'h00}, /* 0x0245 */
            {8'h00}, /* 0x0244 */
            {8'h00}, /* 0x0243 */
            {8'h00}, /* 0x0242 */
            {8'h00}, /* 0x0241 */
            {8'h00}, /* 0x0240 */
            {8'h00}, /* 0x023f */
            {8'h00}, /* 0x023e */
            {8'h00}, /* 0x023d */
            {8'h00}, /* 0x023c */
            {8'h00}, /* 0x023b */
            {8'h00}, /* 0x023a */
            {8'h00}, /* 0x0239 */
            {8'h00}, /* 0x0238 */
            {8'h00}, /* 0x0237 */
            {8'h00}, /* 0x0236 */
            {8'h00}, /* 0x0235 */
            {8'h00}, /* 0x0234 */
            {8'h00}, /* 0x0233 */
            {8'h00}, /* 0x0232 */
            {8'h00}, /* 0x0231 */
            {8'h00}, /* 0x0230 */
            {8'h00}, /* 0x022f */
            {8'h00}, /* 0x022e */
            {8'h00}, /* 0x022d */
            {8'h00}, /* 0x022c */
            {8'h00}, /* 0x022b */
            {8'h00}, /* 0x022a */
            {8'h00}, /* 0x0229 */
            {8'h00}, /* 0x0228 */
            {8'h00}, /* 0x0227 */
            {8'h00}, /* 0x0226 */
            {8'h00}, /* 0x0225 */
            {8'h00}, /* 0x0224 */
            {8'h00}, /* 0x0223 */
            {8'h00}, /* 0x0222 */
            {8'h00}, /* 0x0221 */
            {8'h00}, /* 0x0220 */
            {8'h00}, /* 0x021f */
            {8'h00}, /* 0x021e */
            {8'h00}, /* 0x021d */
            {8'h00}, /* 0x021c */
            {8'h00}, /* 0x021b */
            {8'h00}, /* 0x021a */
            {8'h00}, /* 0x0219 */
            {8'h00}, /* 0x0218 */
            {8'h00}, /* 0x0217 */
            {8'h00}, /* 0x0216 */
            {8'h00}, /* 0x0215 */
            {8'h00}, /* 0x0214 */
            {8'h00}, /* 0x0213 */
            {8'h00}, /* 0x0212 */
            {8'h00}, /* 0x0211 */
            {8'h00}, /* 0x0210 */
            {8'h00}, /* 0x020f */
            {8'h00}, /* 0x020e */
            {8'h00}, /* 0x020d */
            {8'h00}, /* 0x020c */
            {8'h00}, /* 0x020b */
            {8'h00}, /* 0x020a */
            {8'h00}, /* 0x0209 */
            {8'h00}, /* 0x0208 */
            {8'h00}, /* 0x0207 */
            {8'h00}, /* 0x0206 */
            {8'h00}, /* 0x0205 */
            {8'h00}, /* 0x0204 */
            {8'h00}, /* 0x0203 */
            {8'h00}, /* 0x0202 */
            {8'h00}, /* 0x0201 */
            {8'h00}, /* 0x0200 */
            {8'h00}, /* 0x01ff */
            {8'h00}, /* 0x01fe */
            {8'h00}, /* 0x01fd */
            {8'h00}, /* 0x01fc */
            {8'h00}, /* 0x01fb */
            {8'h00}, /* 0x01fa */
            {8'h00}, /* 0x01f9 */
            {8'h00}, /* 0x01f8 */
            {8'h00}, /* 0x01f7 */
            {8'h00}, /* 0x01f6 */
            {8'h00}, /* 0x01f5 */
            {8'h00}, /* 0x01f4 */
            {8'h00}, /* 0x01f3 */
            {8'h00}, /* 0x01f2 */
            {8'h00}, /* 0x01f1 */
            {8'h00}, /* 0x01f0 */
            {8'h00}, /* 0x01ef */
            {8'h00}, /* 0x01ee */
            {8'h00}, /* 0x01ed */
            {8'h00}, /* 0x01ec */
            {8'h00}, /* 0x01eb */
            {8'h00}, /* 0x01ea */
            {8'h00}, /* 0x01e9 */
            {8'h00}, /* 0x01e8 */
            {8'h00}, /* 0x01e7 */
            {8'h00}, /* 0x01e6 */
            {8'h00}, /* 0x01e5 */
            {8'h00}, /* 0x01e4 */
            {8'h00}, /* 0x01e3 */
            {8'h00}, /* 0x01e2 */
            {8'h00}, /* 0x01e1 */
            {8'h00}, /* 0x01e0 */
            {8'h00}, /* 0x01df */
            {8'h00}, /* 0x01de */
            {8'h00}, /* 0x01dd */
            {8'h00}, /* 0x01dc */
            {8'h00}, /* 0x01db */
            {8'h00}, /* 0x01da */
            {8'h00}, /* 0x01d9 */
            {8'h00}, /* 0x01d8 */
            {8'h00}, /* 0x01d7 */
            {8'h00}, /* 0x01d6 */
            {8'h00}, /* 0x01d5 */
            {8'h00}, /* 0x01d4 */
            {8'h00}, /* 0x01d3 */
            {8'h00}, /* 0x01d2 */
            {8'h00}, /* 0x01d1 */
            {8'h00}, /* 0x01d0 */
            {8'h00}, /* 0x01cf */
            {8'h00}, /* 0x01ce */
            {8'h00}, /* 0x01cd */
            {8'h00}, /* 0x01cc */
            {8'h00}, /* 0x01cb */
            {8'h00}, /* 0x01ca */
            {8'h00}, /* 0x01c9 */
            {8'h00}, /* 0x01c8 */
            {8'h00}, /* 0x01c7 */
            {8'h00}, /* 0x01c6 */
            {8'h00}, /* 0x01c5 */
            {8'h00}, /* 0x01c4 */
            {8'h00}, /* 0x01c3 */
            {8'h00}, /* 0x01c2 */
            {8'h00}, /* 0x01c1 */
            {8'h00}, /* 0x01c0 */
            {8'h00}, /* 0x01bf */
            {8'h00}, /* 0x01be */
            {8'h00}, /* 0x01bd */
            {8'h00}, /* 0x01bc */
            {8'h00}, /* 0x01bb */
            {8'h00}, /* 0x01ba */
            {8'h00}, /* 0x01b9 */
            {8'h00}, /* 0x01b8 */
            {8'h00}, /* 0x01b7 */
            {8'h00}, /* 0x01b6 */
            {8'h00}, /* 0x01b5 */
            {8'h00}, /* 0x01b4 */
            {8'h00}, /* 0x01b3 */
            {8'h00}, /* 0x01b2 */
            {8'h00}, /* 0x01b1 */
            {8'h00}, /* 0x01b0 */
            {8'h00}, /* 0x01af */
            {8'h00}, /* 0x01ae */
            {8'h00}, /* 0x01ad */
            {8'h00}, /* 0x01ac */
            {8'h00}, /* 0x01ab */
            {8'h00}, /* 0x01aa */
            {8'h00}, /* 0x01a9 */
            {8'h00}, /* 0x01a8 */
            {8'h00}, /* 0x01a7 */
            {8'h00}, /* 0x01a6 */
            {8'h00}, /* 0x01a5 */
            {8'h00}, /* 0x01a4 */
            {8'h00}, /* 0x01a3 */
            {8'h00}, /* 0x01a2 */
            {8'h00}, /* 0x01a1 */
            {8'h00}, /* 0x01a0 */
            {8'h00}, /* 0x019f */
            {8'h00}, /* 0x019e */
            {8'h00}, /* 0x019d */
            {8'h00}, /* 0x019c */
            {8'h00}, /* 0x019b */
            {8'h00}, /* 0x019a */
            {8'h00}, /* 0x0199 */
            {8'h00}, /* 0x0198 */
            {8'h00}, /* 0x0197 */
            {8'h00}, /* 0x0196 */
            {8'h00}, /* 0x0195 */
            {8'h00}, /* 0x0194 */
            {8'h00}, /* 0x0193 */
            {8'h00}, /* 0x0192 */
            {8'h00}, /* 0x0191 */
            {8'h00}, /* 0x0190 */
            {8'h00}, /* 0x018f */
            {8'h00}, /* 0x018e */
            {8'h00}, /* 0x018d */
            {8'h00}, /* 0x018c */
            {8'h00}, /* 0x018b */
            {8'h00}, /* 0x018a */
            {8'h00}, /* 0x0189 */
            {8'h00}, /* 0x0188 */
            {8'h00}, /* 0x0187 */
            {8'h00}, /* 0x0186 */
            {8'h00}, /* 0x0185 */
            {8'h00}, /* 0x0184 */
            {8'h00}, /* 0x0183 */
            {8'h00}, /* 0x0182 */
            {8'h00}, /* 0x0181 */
            {8'h00}, /* 0x0180 */
            {8'h00}, /* 0x017f */
            {8'h00}, /* 0x017e */
            {8'h00}, /* 0x017d */
            {8'h00}, /* 0x017c */
            {8'h00}, /* 0x017b */
            {8'h00}, /* 0x017a */
            {8'h00}, /* 0x0179 */
            {8'h00}, /* 0x0178 */
            {8'h00}, /* 0x0177 */
            {8'h00}, /* 0x0176 */
            {8'h00}, /* 0x0175 */
            {8'h00}, /* 0x0174 */
            {8'h00}, /* 0x0173 */
            {8'h00}, /* 0x0172 */
            {8'h00}, /* 0x0171 */
            {8'h00}, /* 0x0170 */
            {8'h00}, /* 0x016f */
            {8'h00}, /* 0x016e */
            {8'h00}, /* 0x016d */
            {8'h00}, /* 0x016c */
            {8'h00}, /* 0x016b */
            {8'h00}, /* 0x016a */
            {8'h00}, /* 0x0169 */
            {8'h00}, /* 0x0168 */
            {8'h00}, /* 0x0167 */
            {8'h00}, /* 0x0166 */
            {8'h00}, /* 0x0165 */
            {8'h00}, /* 0x0164 */
            {8'h00}, /* 0x0163 */
            {8'h00}, /* 0x0162 */
            {8'h00}, /* 0x0161 */
            {8'h00}, /* 0x0160 */
            {8'h00}, /* 0x015f */
            {8'h00}, /* 0x015e */
            {8'h00}, /* 0x015d */
            {8'h00}, /* 0x015c */
            {8'h00}, /* 0x015b */
            {8'h00}, /* 0x015a */
            {8'h00}, /* 0x0159 */
            {8'h00}, /* 0x0158 */
            {8'h00}, /* 0x0157 */
            {8'h00}, /* 0x0156 */
            {8'h00}, /* 0x0155 */
            {8'h00}, /* 0x0154 */
            {8'h00}, /* 0x0153 */
            {8'h00}, /* 0x0152 */
            {8'h00}, /* 0x0151 */
            {8'h00}, /* 0x0150 */
            {8'h00}, /* 0x014f */
            {8'h00}, /* 0x014e */
            {8'h00}, /* 0x014d */
            {8'h00}, /* 0x014c */
            {8'h00}, /* 0x014b */
            {8'h00}, /* 0x014a */
            {8'h00}, /* 0x0149 */
            {8'h00}, /* 0x0148 */
            {8'h00}, /* 0x0147 */
            {8'h00}, /* 0x0146 */
            {8'h00}, /* 0x0145 */
            {8'h00}, /* 0x0144 */
            {8'h00}, /* 0x0143 */
            {8'h00}, /* 0x0142 */
            {8'h00}, /* 0x0141 */
            {8'h00}, /* 0x0140 */
            {8'h00}, /* 0x013f */
            {8'h00}, /* 0x013e */
            {8'h00}, /* 0x013d */
            {8'h00}, /* 0x013c */
            {8'h00}, /* 0x013b */
            {8'h00}, /* 0x013a */
            {8'h00}, /* 0x0139 */
            {8'h00}, /* 0x0138 */
            {8'h00}, /* 0x0137 */
            {8'h00}, /* 0x0136 */
            {8'h00}, /* 0x0135 */
            {8'h00}, /* 0x0134 */
            {8'h00}, /* 0x0133 */
            {8'h00}, /* 0x0132 */
            {8'h00}, /* 0x0131 */
            {8'h00}, /* 0x0130 */
            {8'h00}, /* 0x012f */
            {8'h00}, /* 0x012e */
            {8'h00}, /* 0x012d */
            {8'h00}, /* 0x012c */
            {8'h00}, /* 0x012b */
            {8'h00}, /* 0x012a */
            {8'h00}, /* 0x0129 */
            {8'h00}, /* 0x0128 */
            {8'h00}, /* 0x0127 */
            {8'h00}, /* 0x0126 */
            {8'h00}, /* 0x0125 */
            {8'h00}, /* 0x0124 */
            {8'h00}, /* 0x0123 */
            {8'h00}, /* 0x0122 */
            {8'h00}, /* 0x0121 */
            {8'h00}, /* 0x0120 */
            {8'h00}, /* 0x011f */
            {8'h00}, /* 0x011e */
            {8'h00}, /* 0x011d */
            {8'h00}, /* 0x011c */
            {8'h00}, /* 0x011b */
            {8'h00}, /* 0x011a */
            {8'h00}, /* 0x0119 */
            {8'h00}, /* 0x0118 */
            {8'h00}, /* 0x0117 */
            {8'h00}, /* 0x0116 */
            {8'h00}, /* 0x0115 */
            {8'h00}, /* 0x0114 */
            {8'h00}, /* 0x0113 */
            {8'h00}, /* 0x0112 */
            {8'h00}, /* 0x0111 */
            {8'h00}, /* 0x0110 */
            {8'h00}, /* 0x010f */
            {8'h00}, /* 0x010e */
            {8'h00}, /* 0x010d */
            {8'h00}, /* 0x010c */
            {8'h00}, /* 0x010b */
            {8'h00}, /* 0x010a */
            {8'h00}, /* 0x0109 */
            {8'h00}, /* 0x0108 */
            {8'h00}, /* 0x0107 */
            {8'h00}, /* 0x0106 */
            {8'h00}, /* 0x0105 */
            {8'h00}, /* 0x0104 */
            {8'h00}, /* 0x0103 */
            {8'h00}, /* 0x0102 */
            {8'h00}, /* 0x0101 */
            {8'h00}, /* 0x0100 */
            {8'h00}, /* 0x00ff */
            {8'h00}, /* 0x00fe */
            {8'h00}, /* 0x00fd */
            {8'h00}, /* 0x00fc */
            {8'h00}, /* 0x00fb */
            {8'h00}, /* 0x00fa */
            {8'h00}, /* 0x00f9 */
            {8'h00}, /* 0x00f8 */
            {8'h00}, /* 0x00f7 */
            {8'h00}, /* 0x00f6 */
            {8'h00}, /* 0x00f5 */
            {8'h00}, /* 0x00f4 */
            {8'h00}, /* 0x00f3 */
            {8'h00}, /* 0x00f2 */
            {8'h00}, /* 0x00f1 */
            {8'h00}, /* 0x00f0 */
            {8'h00}, /* 0x00ef */
            {8'h00}, /* 0x00ee */
            {8'h00}, /* 0x00ed */
            {8'h00}, /* 0x00ec */
            {8'h00}, /* 0x00eb */
            {8'h00}, /* 0x00ea */
            {8'h00}, /* 0x00e9 */
            {8'h00}, /* 0x00e8 */
            {8'h00}, /* 0x00e7 */
            {8'h00}, /* 0x00e6 */
            {8'h00}, /* 0x00e5 */
            {8'h00}, /* 0x00e4 */
            {8'h00}, /* 0x00e3 */
            {8'h00}, /* 0x00e2 */
            {8'h00}, /* 0x00e1 */
            {8'h00}, /* 0x00e0 */
            {8'h00}, /* 0x00df */
            {8'h00}, /* 0x00de */
            {8'h00}, /* 0x00dd */
            {8'h00}, /* 0x00dc */
            {8'h00}, /* 0x00db */
            {8'h00}, /* 0x00da */
            {8'h00}, /* 0x00d9 */
            {8'h00}, /* 0x00d8 */
            {8'h00}, /* 0x00d7 */
            {8'h00}, /* 0x00d6 */
            {8'h00}, /* 0x00d5 */
            {8'h00}, /* 0x00d4 */
            {8'h00}, /* 0x00d3 */
            {8'h00}, /* 0x00d2 */
            {8'h00}, /* 0x00d1 */
            {8'h00}, /* 0x00d0 */
            {8'h00}, /* 0x00cf */
            {8'h00}, /* 0x00ce */
            {8'h00}, /* 0x00cd */
            {8'h00}, /* 0x00cc */
            {8'h00}, /* 0x00cb */
            {8'h00}, /* 0x00ca */
            {8'h00}, /* 0x00c9 */
            {8'h00}, /* 0x00c8 */
            {8'h00}, /* 0x00c7 */
            {8'h00}, /* 0x00c6 */
            {8'h00}, /* 0x00c5 */
            {8'h00}, /* 0x00c4 */
            {8'h00}, /* 0x00c3 */
            {8'h00}, /* 0x00c2 */
            {8'h00}, /* 0x00c1 */
            {8'h00}, /* 0x00c0 */
            {8'h00}, /* 0x00bf */
            {8'h00}, /* 0x00be */
            {8'h00}, /* 0x00bd */
            {8'h00}, /* 0x00bc */
            {8'h00}, /* 0x00bb */
            {8'h00}, /* 0x00ba */
            {8'h00}, /* 0x00b9 */
            {8'h00}, /* 0x00b8 */
            {8'h00}, /* 0x00b7 */
            {8'h00}, /* 0x00b6 */
            {8'h00}, /* 0x00b5 */
            {8'h00}, /* 0x00b4 */
            {8'h00}, /* 0x00b3 */
            {8'h00}, /* 0x00b2 */
            {8'h00}, /* 0x00b1 */
            {8'h00}, /* 0x00b0 */
            {8'h00}, /* 0x00af */
            {8'h00}, /* 0x00ae */
            {8'h00}, /* 0x00ad */
            {8'h00}, /* 0x00ac */
            {8'h00}, /* 0x00ab */
            {8'h00}, /* 0x00aa */
            {8'h00}, /* 0x00a9 */
            {8'h00}, /* 0x00a8 */
            {8'h00}, /* 0x00a7 */
            {8'h00}, /* 0x00a6 */
            {8'h00}, /* 0x00a5 */
            {8'h00}, /* 0x00a4 */
            {8'h00}, /* 0x00a3 */
            {8'h00}, /* 0x00a2 */
            {8'h00}, /* 0x00a1 */
            {8'h00}, /* 0x00a0 */
            {8'h00}, /* 0x009f */
            {8'h00}, /* 0x009e */
            {8'h00}, /* 0x009d */
            {8'h00}, /* 0x009c */
            {8'h00}, /* 0x009b */
            {8'h00}, /* 0x009a */
            {8'h00}, /* 0x0099 */
            {8'h00}, /* 0x0098 */
            {8'h00}, /* 0x0097 */
            {8'h00}, /* 0x0096 */
            {8'h00}, /* 0x0095 */
            {8'h00}, /* 0x0094 */
            {8'h00}, /* 0x0093 */
            {8'h00}, /* 0x0092 */
            {8'h00}, /* 0x0091 */
            {8'h00}, /* 0x0090 */
            {8'h00}, /* 0x008f */
            {8'h00}, /* 0x008e */
            {8'h00}, /* 0x008d */
            {8'h00}, /* 0x008c */
            {8'h00}, /* 0x008b */
            {8'h00}, /* 0x008a */
            {8'h00}, /* 0x0089 */
            {8'h00}, /* 0x0088 */
            {8'h00}, /* 0x0087 */
            {8'h00}, /* 0x0086 */
            {8'h00}, /* 0x0085 */
            {8'h00}, /* 0x0084 */
            {8'h00}, /* 0x0083 */
            {8'h00}, /* 0x0082 */
            {8'h00}, /* 0x0081 */
            {8'h00}, /* 0x0080 */
            {8'h00}, /* 0x007f */
            {8'h00}, /* 0x007e */
            {8'h00}, /* 0x007d */
            {8'h00}, /* 0x007c */
            {8'h00}, /* 0x007b */
            {8'h00}, /* 0x007a */
            {8'h00}, /* 0x0079 */
            {8'h00}, /* 0x0078 */
            {8'h00}, /* 0x0077 */
            {8'h00}, /* 0x0076 */
            {8'h00}, /* 0x0075 */
            {8'h00}, /* 0x0074 */
            {8'h00}, /* 0x0073 */
            {8'h00}, /* 0x0072 */
            {8'h00}, /* 0x0071 */
            {8'h00}, /* 0x0070 */
            {8'h00}, /* 0x006f */
            {8'h00}, /* 0x006e */
            {8'h00}, /* 0x006d */
            {8'h00}, /* 0x006c */
            {8'h00}, /* 0x006b */
            {8'h00}, /* 0x006a */
            {8'h00}, /* 0x0069 */
            {8'h00}, /* 0x0068 */
            {8'h00}, /* 0x0067 */
            {8'h00}, /* 0x0066 */
            {8'h00}, /* 0x0065 */
            {8'h00}, /* 0x0064 */
            {8'h00}, /* 0x0063 */
            {8'h00}, /* 0x0062 */
            {8'h00}, /* 0x0061 */
            {8'h00}, /* 0x0060 */
            {8'h00}, /* 0x005f */
            {8'h00}, /* 0x005e */
            {8'h00}, /* 0x005d */
            {8'h00}, /* 0x005c */
            {8'h00}, /* 0x005b */
            {8'h00}, /* 0x005a */
            {8'h00}, /* 0x0059 */
            {8'h00}, /* 0x0058 */
            {8'h00}, /* 0x0057 */
            {8'h00}, /* 0x0056 */
            {8'h00}, /* 0x0055 */
            {8'h00}, /* 0x0054 */
            {8'h00}, /* 0x0053 */
            {8'h00}, /* 0x0052 */
            {8'h00}, /* 0x0051 */
            {8'h00}, /* 0x0050 */
            {8'h00}, /* 0x004f */
            {8'h00}, /* 0x004e */
            {8'h00}, /* 0x004d */
            {8'h00}, /* 0x004c */
            {8'h00}, /* 0x004b */
            {8'h00}, /* 0x004a */
            {8'h00}, /* 0x0049 */
            {8'h00}, /* 0x0048 */
            {8'h00}, /* 0x0047 */
            {8'h00}, /* 0x0046 */
            {8'h00}, /* 0x0045 */
            {8'h00}, /* 0x0044 */
            {8'h00}, /* 0x0043 */
            {8'h00}, /* 0x0042 */
            {8'h00}, /* 0x0041 */
            {8'h00}, /* 0x0040 */
            {8'h00}, /* 0x003f */
            {8'h00}, /* 0x003e */
            {8'h00}, /* 0x003d */
            {8'h00}, /* 0x003c */
            {8'h00}, /* 0x003b */
            {8'h00}, /* 0x003a */
            {8'h00}, /* 0x0039 */
            {8'h00}, /* 0x0038 */
            {8'h00}, /* 0x0037 */
            {8'h00}, /* 0x0036 */
            {8'h00}, /* 0x0035 */
            {8'h00}, /* 0x0034 */
            {8'hfd}, /* 0x0033 */
            {8'h1f}, /* 0x0032 */
            {8'hf0}, /* 0x0031 */
            {8'h6f}, /* 0x0030 */
            {8'h00}, /* 0x002f */
            {8'h02}, /* 0x002e */
            {8'h80}, /* 0x002d */
            {8'he7}, /* 0x002c */
            {8'h00}, /* 0x002b */
            {8'h02}, /* 0x002a */
            {8'ha2}, /* 0x0029 */
            {8'h83}, /* 0x0028 */
            {8'h18}, /* 0x0027 */
            {8'h80}, /* 0x0026 */
            {8'h02}, /* 0x0025 */
            {8'h93}, /* 0x0024 */
            {8'h10}, /* 0x0023 */
            {8'h50}, /* 0x0022 */
            {8'h00}, /* 0x0021 */
            {8'h73}, /* 0x0020 */
            {8'h30}, /* 0x001f */
            {8'h42}, /* 0x001e */
            {8'h90}, /* 0x001d */
            {8'h73}, /* 0x001c */
            {8'h00}, /* 0x001b */
            {8'h82}, /* 0x001a */
            {8'h82}, /* 0x0019 */
            {8'h93}, /* 0x0018 */
            {8'h00}, /* 0x0017 */
            {8'h08}, /* 0x0016 */
            {8'h02}, /* 0x0015 */
            {8'hb7}, /* 0x0014 */
            {8'h30}, /* 0x0013 */
            {8'h04}, /* 0x0012 */
            {8'h60}, /* 0x0011 */
            {8'h73}, /* 0x0010 */
            {8'h30}, /* 0x000f */
            {8'h52}, /* 0x000e */
            {8'h90}, /* 0x000d */
            {8'h73}, /* 0x000c */
            {8'h02}, /* 0x000b */
            {8'h02}, /* 0x000a */
            {8'h82}, /* 0x0009 */
            {8'h93}, /* 0x0008 */
            {8'h00}, /* 0x0007 */
            {8'h00}, /* 0x0006 */
            {8'h02}, /* 0x0005 */
            {8'h97}, /* 0x0004 */
            {8'hf1}, /* 0x0003 */
            {8'h40}, /* 0x0002 */
            {8'h25}, /* 0x0001 */
            {8'h73}  /* 0x0000 */
        };
        
        localparam int unsigned NumBytes = DataWidth/8;
        localparam int unsigned WordOffset = $clog2(NumBytes);
        logic [BootromSize/NumBytes-1:0][DataWidth-1:0] rom_word_addressed;
        assign rom_word_addressed = rom;

        logic [$clog2(BootromSize)-2:WordOffset] aligned_address; // Bootrom is only half size.

        assign aligned_address = addr_i[$clog2(BootromSize)-1:WordOffset];

        assign data_o = rom_word_addressed[aligned_address];
        
    endmodule
