`ifndef CSR_DEF_SVH
`define CSR_DEF_SVH

`define Address_A_CSR 32'h3c0
`define Address_B_CSR 32'h3c1
`define Address_C_CSR 32'h3c2
`define B_M_K_N_CSR 32'h3c3

`endif