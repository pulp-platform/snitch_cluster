`ifndef CSR_DEF_SVH
`define CSR_DEF_SVH

`define Address_A_CSR 32'h3c0
`define Address_B_CSR 32'h3c1
`define Address_C_CSR 32'h3c2

`define B_M_K_N_CSR 32'h3c3

`define ldA_CSR 32'h3c4
`define ldB_CSR 32'h3c5
`define ldC_CSR 32'h3c6

`define StrideA_CSR 32'h3c7
`define StrideB_CSR 32'h3c8
`define StrideC_CSR 32'h3c9

`define STATE_CSR 32'h3d0

`endif